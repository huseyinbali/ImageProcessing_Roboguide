��  	c4�A��*SYST�EM*��V9.1�0214 8/�21/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP6fBI�IZ@!�LRM_RECO�"  � ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� ."��!_I�F� � 
$_ENABL@C#T� P dC#U5K�!CMA�B �"�
� �OG�f 0CUR�R_D1P $Q3LI�N@S1I4$C$AU�SOd�APPI�NFOEQ/ 9�L A ?1�5�/ H �7�9EQUIP �2�0NAM� ���2_OVR�?$VERSI� �� PCOUPLE�,   $�!PPV1CES C G�1�!�PR0�2	� � $SOF�T�T_IDBTOTAL_EQ� �Q1]@NO`BU SPI_INDE]�uEXBSCREE�N_�4BSIG��0O%KW@PK�_FI0	$�THKY�GPAN�EhD � DUMMY1d�D�!U�4 Q!RG1R�
� � $TIT1d ��� 7Td7TP� 7TP7T55V65VU75V85V95W05W�>W�A7URWQ7UfW1*pW1zW1�W1�W �6P!SBN_CF��!�0$!J� ; 
2�1_CMN�T�$FLAG�S]�CHE"�$Nb_OPT�2p��(CELLSE�TUP  `f�0HO�0 PRZ1}%{cMACRO�bOREPR�hD0D+`t@��b{�eHM �MN�B
1�UT�OB U��0 9DEVIMC4STI�0�� �P@13��`BQdf"V�AL�#ISP_UsNI�#p_DOv<7IyFR_F�@K%�D13�;A�c�C_�WA?t�a�zOFFu_@N�DEL�x�LF0q�A�qr?1q�p�C?�`�Ab�E�C#�s�ATB�t��d�MO� �sE' � [M�s���2�REV�BI�LF��1XI� %�R�  � OD�}`j�$NO`M�+��b�x�/�"u�� ����!�X�@Dd p =E RD_Eb��?$FSSB�&W`�KBD_SE2uAUG� G�2 "_��B�� V�t:5`ׁ�QC ��a_ED|u � � C2���`S�p�4%$<l �t$OP�@QB9�qy�_OK���0, P_C� y��dh��U �`LACI�!��a���� FqCOM9M� �0$D��ϑ��@�pX��OR BI�GALLOW�� (KD2�2�@V�AR5�d!�AB e`BqL[@S � ,K�JqM�H`S�pZ@M_�O]z���CFnd X�0GR@���M�NFLIx���;@UIRE�x84�"� SWIT=$�/0_No`S�"CFzd0M� �#PEED��!�%`(���p3`J3tV�&$�E�..p`L��ELBOF� �m�� m�p/0��CP�� F�B����1��r@1oJ1E_y_T>!�Բ�`��g���G�� �0WARNMxp�d�%`�V`wNST� COR-�rFLTR�T�RAT T�`� $ACCqM�� R�>r$ORI�.&�ӧRT�SFg�_��CHGV0I�Ep�T��PA�I{��T�!��� �� �#@a���HSDR�B��2�BJ; ��C��3�4�5��6�7�8�9�>���x@�2 @.� TRQ��$%f��4ր����_U����z��Oc <� �����Ȩ3�2��LL�ECM�-�MULTIV4�"$��A
2q�CHILD>�
1���z@T_1b  4� STY2�b4�=@�)24����@��� |9$��T��A�I`�E��eTOt���E��EXT����ᗑ�B��22(�0>��@��1b�.'��B ��A�K�  �"K�/%�a��R� ��?s!>�O�!M��;A�֗�M�� 	� � =�I�" L@�0[�� R�pA��$JOBB�����`�v��IGI�# dӀ ����R�-'r��A��ҧ��_M��b$ �tӀFL6�BNG�A��TBA� ϑ� !��
/1�À�0����R0�P/p ����%�|��Bq@W��
2JW�_RH�C�ZJZ�_zJ?�D/5C�	�ӧ��@�����Rd&� �����ǯ�rGӨg@N�HANC��$LG /��a2qӐ� ـ@��!A�p� ���aR��0>$x��?#DB�?#3RA�c?#AZt@�(p.�����`FCT��ƕ�_F࠳`�SM��!I�+lA�%` � ` ���$/�/����[�a��M�0\��`l��أHK��AEs@�͐�!�"W��N� S�'�I��'  E. II��2�(p�STD_C�t�1Q���USTڒU�)�#�0U[�%?IO1��� _Up�q��* \��=�AOR@zsBp;�]��`O6  RSY�G�0�q>E�Up��H`G�� {@]�DBPXWORK��+��$SKP_l�p��DB�TR�p , �=�`����Z m�OD3��a �_C"�;b�C� �GPAL:c�a�tőS�D��G�Bb����Pl�.� )DB�!��-|B APR��
p�@Ja3��. /��u����� �LUY/�b_tS��0�_����PC�1�_�TEsNEG�]� 2�_̹S6PRE.��R3�H $C��.$Lc/$USނz �)kINE�7A_D1%�ROyp��������qbc7 T@zfPA����RETURN\xb�MMR"U��vI�CRG`EWM�0^�SIGNZ�A ����e� 0$=P'�1$P� m�2�`��`tm�pDIp �'�Bd.a	r>�GO_AW ����0ؑB1m@CS,d�(�CYI�4���`�1wsqu�|t2vz2��vN�}��E]sD�EVIS` 5 oP $��RB���I�wPk��vI_#BY���p�TQ�t�HNDG�Q6 �H4��1�w��$DSBLC��O��vG@h�Ǝ@_qL��7/��F@]�d�FB���FERa8����t]s����8> i�T1?���MCS솀�FD ���[2H� W��EE���%8F��ŻtSLAd��0w9  ��INP^���]�`�]q��:P +8�S��0x�^���^���FI�2��������A	AW�l���NTV�㜒V�~���SKI�#TE�����a���T1J_�#;2_�PD�SAF��T�_SV�EX�CLU�῰�D6@Ll �Yք��3��HI_V
0\2PPLY�@0«�G������_ML%��pVR�FY_�C��M��I3OC�UC_� �d��O�p��LS�`�V�&T4�A1��s����@PdE&�gp�AU��NFT�u��uZ�8�pm�ACHD�O�؆�^���AFC CPl��TD�4P~�� ��' ;�P@T�ѡ0�,@ ���}�N���=� <Y���TĲ�?� ���{�SG5N��=;
$�` �a>aR0I�3�g@ _B�M�_B]�ANNUN��P~��ÅuC.@ �`/�ɢ�� �����2�EFC@I�R>p�c$F���4OT�`�{�&TD�(RQ<�#QdZJ�Mb�NI�R?���4һ6�A��R�DA=YCLOAD�tT�-�'S5#Q�EF_F_AXI��@�P�QO3O�йS�@_�RTRQ��A D�1�	`��Q,@ B��EVp�Ӓ���@�0`}�0��{��MP�E{� BV����0�$s��DU�`��]��BCAB��C��f�PNS"�+0ID�CWR���V!� V�w�V_���V �DI�� �4D� 1$-V�`SEm�TQ�j}�'���D�^E�_n�$�VE� � SW���[a�d����A��OH��f)�PP��%�IR�1Bu@p�&���b�� ��]�w3W�O � W��v�M���C�0��cp��R7QDWF�MSw0���AX,���$�LIFAE�@����-Q��N�� ����Co���-CB0LqN]a̐��OV0HE�Q�SUP�T�D���@_oS�1_�(�Gq�Z�
W�
B1`��#��@�k2XZ_ �LQY2�C9`T�_@``��N�����J
�! >�_� ��F� ބ4E `�pCA�CH,�\�]SIZ�(T ���bN�UFFI� ���@(HT��'S6#Q�BMp0��F 8��KEYoIMAG�cTM,a�V#��a�^�hB1�OOCVIE�aG�2� L��H���?� �	��D� PH��6�ST'�!C"D��K$PK$-�K$��K EMAILK�u`[��0^��FAUL�RI�28sc�C� COU�0iA��0T`�1J< �$�#�S�m�ITW�BUFp��p(�t�0�0n B�$�t�C�����"�3� SAV-5�"����H7@@��P44�
`�N�a_� 5LЉ9OTgb+���P�P�:���7#AXC����X� T��a3_G��
m@YN�_N� K <\�D��uPb�M�M8�jH TL�F~`$�`��DIزE�@`��aLY���G1��&�G�Da:AF����baM��`A�#�3C_^`�`Knd�@^DQ��R��E�(ADSPl�BPC�KIM:3 �C�A��A��U�Gd meڠ� IP��C7�3�DTH���B�ЙTaa�CHSEC�CB#SC	�"�PV���Z`�P�3�Tp��NVk�AG�S�T�F� F����0d�C5@�1aSC8���u�CMER��Q�FBCMP��~@E�T;� N�FU� DU� ́�`����CD�IYP�0�#d���`NOu�=�O�� �pzbL�xds�P�zbEC"��e
��2�!�uc�0� PH *�aL��_c�q�1f�� ,�'��dD��f"��f-Ѡ�f���f��f7�i8B�i9�j���hz1zU1z1(z15z1BzU1Oz1\z1iz2wz�2{z2z2(z2�5z2Bz2Oz2\z2*iz3wz3z3{zU3(z35z3Bz3Oz�3\z3iz4wr�EXT��=�QB\h@@%@�e@C��e�0�FDR��RT� VW��2�򁑇R��REM��Fq��O�VM�C��A��TR�OV��DT80КMXߜIN��: Ϛ��'IND���
�F@�0@G�1d�ِ9 r��D��ِRIV԰�&��GEAR�AI%O��K��$�N5@���������� %�Z_�MCM� ���Fve UR3bS ,�a�1? 9 P?����?�E@,����1`v�T�j��P�1��RI^e����#ETUP2_� U -��#TDGP0��$Ti��Z�T��qa�"BACBV QTD��"eD)_J%��8�c0@ѰIFI:�0@0`�`�Ь�PT���LUI6$W �� (� URt�1@@�2MA�P� ����I��u$(�Sܰ?x4��Jb@CO|0�3VR�T$���x$SHO8�ѱ��#ASSjP�18(IPQ�BG_�����s��s��(s��5sF�ORC�"7��DAkTA��X�"FUס�1:B��2:ALOG����Y |*�N;AV�0�(�X�����S�"&$VgISI[�.BSC�4�SE�t�7�VB�O
r���Bò�A�Z֯$PO,�IE���FMR2s�Z ��i`f⁑ s@�օ�������ǖ� ��堒_wqX���I#T_ֱSd��ME�j��|�DGCLF;�D7GDYd�LD�H�!5
?�ѡMcp8#�[��� T�sFS�07$\ P2����sC�0$EX_������1�0�PE��53�5��G�Q��g] ��0bSW5}O��DEBUG��L]�GRc��U�S�BKU`O1�p  PO�Ј�t��"`G�t�Ms�LOO,�3��SM�E<2|���& _E ^ y��TERM��9_��� ORISA��y`��cp�SM_`@�]���a������ b���~�UP"c�3 -�D�^(����f _>�Gk
}�EL�TO�!>B�PFIGf?AנS�`b�`$UFRfB�${`�� Ne�OT���PTAiP���N;STT@PAT^Qi��PTHJ&aL`Ep9 d2U`�ARTU0��� U1�">AREL<Ac1SHFTPR?A3__�R/`Ic% ) $8�b.႐8S�S�2SHId+��U�b O1AYLO .P�1 A��j����e[PERV p�� �$��T@A��Ȱ+%̫�ȰRC��eAScYM3A�e?AWJ�$� �E$�/[)�OaU$T@ A3��&IaPS��Q�ORT@�M��/����d���t��� �16�H9Os���e �˶,s�i`OC���$OP^��A�cFv���a�i@��2R0R�S"OU�Se�R�5m8K���e$PWR]�IM�5"R_H3(*И ?AUD$�kS�Voc1SDfH�$�HdE!@ADDR
C�H��G7A,A%Ap"�p@F��ag H2�S�PFѝ�dE��dEs�dE(sSE��H��`H�SY`MN�h�W�@0��"QebaOL�/SW�{0R�\f��AC�RO����ND_�C/Szb��4�QROUP�S2_��
Ғ�11�q��:S�DY3  DY��EXpDY(pDY��⊒AC���SAVE�D?W�SOUG�C��gi $��@0_D)�x��j«BPRM_
�}~�HTTP_z`�H�aj (;`OB�JB�%B��$C�L�E�0a�`k �� 4��6�_�TĽ�XbS0�3��KR�L�9HITCOU����G�LS�j0Xbb�`$�f�j0ʷk0SS����dJQUERY_�FLA�C_ _WE�BSOCI��HW�cq�+�l_@� IONCPU�R*�Ov ma��K�0pzD/q�D/q~ǂ�IOLN���m 82�R��i��$SL��$INoPUT_��$�0�~xPy� dZpS)L�P+�nep{�u`�tB#�uB"NAIO�P�F_AS��o��Q$��B��qN�Yр�2��ksM�ts�H�YB�5���A�pUOP��p `�pS�C�@��%���,�}��0P�3��0s���,������I�P_ME\��q �X�pIP,@�Rւ_!NP��`*�G2B��O��BSP���P��F�BG�Q�-�M<!��r l �TA4�3`As�TI���%�� ��_�OPS^�BU��ID�Ўbs����x0��;a-���� sD�r?�r�S��pNҘ���ӕ�IRCA_�CN� t ��Ji�pCY�@EA ��C��q��31�#���@z"���!DAY_<����NTVA�����u��r#��u�SCA��u�CLO᎑j����@��u��ڔ$��N_R0Cβ򐎒c�6�v�r��^3%����'b�����Pi��� 2u �p.�����w��\�'b\�LABp�z��Ѐ�UNIб9n�	 ITYl�.�D0EL�R; G���x�r��R_URLЀ$A�AEN|�k�*�t�0�CT�AT_U#§ �Jp��yр!$�_%E�pRk�.�"�AS��q8�J�aC�#FL��K��P
W�r��
�UJR�%z �J`F��(����=D£$J7S%�J8��7&�h������7���8�ɭ�AP�HI�Q����D���J7J8"�L�_KE��  ��KQpLMܑ 7{ <٠XR�p$p��WATCH_V�A�A�ű#fFIE�L�"Cy�2Ҳ�|� 
��V�G-1��C�Tܰ������LG~ɳ}� !�?LG_SIZRdv�`�հ����p��FD��I���ة��������� ��d3��V��V��pV��V���V�K!G�� _� _CM�����ꂫ�F�!�����А4(�Ѡ������ ���p��� �I��
�`����������RSU��  (��LNԢ��"~_��`DE��E�r!�s���S��r0L���DAU���EA�PQp44���GqH52X��pBOOYA?� C�ʀ�IT�c��� �RE4�SCR��|c��D�PKr,QMARGI�q�;�v�S4e$�d�qS8c�rWC�qܕ��JGM�MN3CH���qFN(Ҟ1K����	UF��n�FWD�HLSTP�
V����,���RS?H� ��C�~"�� w�U�Q�v���d��G�	PPO��"2�� ��	E]X�TUI�I;� ��;�8bZ#�Z#� ���R��P# #9N�A�3ANA�rA1���AI���D�� �D�CSf�lC�#zC�"O��(O�'SK�2�(S�(ZIGN�Ў��0���4��$DEA|�LL"�Xp�q���Ѐ4�м�T��$�׳��r
���AA�B��۠lp*s�A��+S1�52�53�1.�8"� �Ђ �Jk�0�$�u�t���Q�e����:FSTe�R��Y�B\A �$EkFCkK���PzFp�F{�$�у Lp #�n�8����Co`��d��P�D�5#_ ��X�Np�Q��$ So��MCt�� ��J`CLDPe� �TRQLI��"�PY>T�FL%�iR�QrS��D��rWpLDrU\TrU�ORG(�v�R��RESERV2t�T>s��TIr /Sv�� �� 	[UvMTrUS�Vd�PP^�	�Q+d>3fRCLMCAd�_��_SiTp3al0MDB�G�qͰ�?�$DEBUGMAS&�(_�P���UuT� |��E����PFRQ~V�� � �ٿHRS_RU�q��A'�A5��FRE�Q����$� ��OVERt���F���P�EFI��%��A(��a�T�a�T� q\�q��$U@�%�?`��PS�0C�	sC��BcN��sScUݐ�a?({ 	�1MISCu�g� d}�ARQA��	�TBN �� �m!�AX �-��>.�EXCES�{�R�rM��̱����r� Ŀ��rSC@ '� H"�	�_S���8���,�>�.PKɴ���r��N �eB_��F�LIC�DB QU�IRE�MO��O��pv�QL�@Mȵ� P��E����Ab��aND��q�ހ��{�r��؄�D���I�NAUT4��RSM����+0N$bn�xj�|�r�PSTḺw� 4٠LOCF�RI��EEX�A�NG�"�q�aODA�e��p|����MF���Cv7I�BA p�Eq�o�fSUP�Fv?�FX;�IGG � �`�Cn� (�C��Da�br\B�� ^@ɨ^@ئ���P��7��qTIvл�[�o�M�+��b� t9�MD6���)D�� O�XaL�qH���O�DIA��P�>�WiO��1�O�D��)|�Ot�)`ހ�� m�CU��V ��#`�q��\_�`y�� ���CC��`rr�� �P �J���P��KE�^����-$B+p��@ND�2ZbZ�P�2_TX�DXTRA�#|�lbM�E�LO��ހ�k�$�����u�ǲ��ܪ�ߒRR2�u��� .����A0a d$CALI��o�G�!��2�0RI�N����<$R��S�W0_d,�lcABCJ�D_Jb����pC��_J3W�
Q�1S�P�Т��pPQ�x�3Pw�̱�@�p��Jlch���R(aOu1IMl`�rCSKP_Z�Ի�$�#��J���rQ���p�����_AZ/b���I�ELZ1��ZaO�CMP��q�q��R1T�at��1��В�F�1���{ ��Z���SMGY'�zdJG�PSCLN�
�SPH_0�p7��㓰�p=��RTER+���I� ��_� )Q6@aA\ SC�r'�DI_�n��23U��DF�0�H�LWN�VEL�PQIN�Bf q�_BAL� �ry��ѳqJi�x~�����MECH�2?�N�IN
�q��!�ǲ��]�q��@_�p �����/���@�􆂛��?���D�HN�~�����0$aV������{!$��X'qrA�$O1����u�H �$B�ELZ��g�_ACCE� �la� OIRC_(��a�P�NT�q;C$PSN�CRL�0��XS ���?�� �G��	D�3�ؠQ�_�1�lIO"u�p�_M�GsDDl(�rFW3P(�����}�DE�PPABN6�RO��EE_�1 �PP��1�a����0?$USE_���#]P+pCTR�$Y��~ .a �AYN�pA m 6&��f�6!M�aұ��"fOk�
c$INC�������'��.�ENC�L��r����� INCBI0��%)���NTi��NT23_L�r�#CLO]�r09pI\� �6R���p���0���C���&MOSI�q��߰O!s�rPERCH  ��7q� y7��3�2zd�@o�g� %&N��AC�5L$�ӻ����%��8:F36TRK��AAY���3��HACWE�LC�z暁�"�`MOM}"����P̰�����cC���DU���DS_BCKLSH_CC�E�`X6 8p>#�s�C�"ZM!�CLALM�$�a�@ 5UCHK���Z�GLRTY��A��$���Q'�_f�M4_U	M�c�VC�cz��SnpLMTt�_Lj b�Tv��WE�]�P�[ �P��U��нc�2 d&�8PC�1�8H��&�p�UCMC��z~CN_	�N��f��SF��9V "��'��TaC�eXhCAT�^SHf�	�~�&yQ��A�&����ɗ�mP�A�T�"_P�UrC_ ����OFm0��_CqtbU�JGJ�d�esW�OG|rg�TORQU  ��K3hI��c2��r_W�EHD��m�tP^�ud�uI�{I
�IdF0��q��I���vVC� 0����j��1p�n��0�v�JRaKp�������DB���M����M��_DL^�2GRV�t�^�dՁH_��Ӄ�"�COS/�|�/�LN��R�s�Y�^ T���@T�&���~�D�ЅZM�c6ՁMY[�Θ;�I�|C��THET0#5NK23d�X\�[CB�CBXC��AS�C�&�Q�^Q���SB^o�)�GT	S���C{�Kq��:sx�祪��$DU_P@�7ʢ��٧��Q�1Y_4cqNE��AKoT��-�< �A��:�C�!�,�,�LPH/���%�Ss���~� �������������:�EV\�VQ�N t�V��UV��V��V��V��VȻVֹH\�u�{�Ps��a�Ȑ�H��H��UH��HȻHֹOM��O\�O�r�O��O���O��O��O��O
ȻO��F�>���~����O�SPBALA�NCE_ޑ��LE6��H_�SP��o����~��ҍ�PFUL�C����⍕��1=���UTO_ZPbU�T1T2^�2N AQ�� ~���A���(���AT	@OA�>�pINSEG�<1�REV��<0�!DI�F2E	1���?�1�%@OB��%Q���G�2�p� LQ݄LCHgWAR�SABAq�E��<0ސU!����XUAPdt�3�?S��� 
u��q��%ROBm0CRC��ib�VP�C�_]rT �� x $W�EIGHR p$�M���tpIR!0IF�
!�LAGC""bS�C"��C"BIL)O1D�@?0ST� P��%P {�`��������
� �D!]q � 2�J4DEB�ULXɠM'MY9���N+s��p$D�1$�� op � ��D�O_� A�� <@��rh��D!0�BB�: N�#_!0D 3�_O2P ��� %�PT� �!�QTx��� TICK-�T1� %j�@s!Nm0M�	m0R�@D!�=�=�� PRO�MPR#E/� $IR�pB!hP��0"MAIڀ}!T"�_# ���^AV �R�CODwFUJ ID_�0'%������G_SUFF�&� 9!��DO����< �GR#=�e$�q$=�|%=�%�qe$�� ����H�_FIv�9�#ORDB ��36b�"B!� $ZDT.%�_���4 *��L�_NAs52�DEF_IE852�Q4 �I�S�}3��5�IS��`��D�3�O4�a�4�a�bSDQ��B�4wD�pO�� LOCKE+q_#����1e"_ UMd%52e$}3e$ �5e$�2q"gCp%`3q$ �4q"Q�F�1|#H�^q |%52|%}3|#�GUa(8P�4H�1�� �WFHEU<Cxp�T�E0Q�� >LOMB__RzW�0VIS=�IT�YAoqOCA_�FRIN�S�SI�1�Q�Rp�W{�W)3�W�XW�[��V��_i�!EAS �"�q�Tp@��V�4�Y5�Y6OR�MULA_I+q��G%7� h ��7�COEFF�_OW��dW��GdqS �CA����_GR� ?� � $<@��
XGTM/G't<E�]DCA|ER��T�%D$4� �  G�L�L�$@S/�_SVL�4�x$hV� �ܒd� � rSE;TU�3MEA�D �b� _�"�� �3 �p�� � �`@ �� �A�:2s$A0AD�b�Q�";��@�1@G��:��REC�!�=��MSK_��s�� P��1_USERz�j���,���z�VEL>���,������=�I0f��M�T8CFG��� � u��Oc�NGORE�� ��-�~�� 4 �s8^�d�XYZ�#f����d� �_ERR�� ��ep6 A�c\�}��Ҁ� BUFINDX1����W�MORt� H��CU\�d�����1Ӄ���!$���10��a���Gr� � $SI�`�P ��Ɲ�VO
����OB�JE��ADJU���AY9p���DJ�OU� 5���C!.�"=��T��y�8��x��DIR}���p�������DYNb$�b��TR�5�R�QH�B 4��OPWOR�� �,� S�YSBU*�2�SO!P���q�U���1P<@߂4�PA���X6�_�2�OPz U4��(��t�e�IM�AGo���q�SIM��IN`\���?RGOVRD��%���g�Pi��������@( C׵d�L:@BY���> �PMC_E0���N*�M±�1���p��SL����{ ���OVSL��S:RDEX�1�0K�2c���a_��cǬ  ��cì mÂ�}Ȫ�ÁC��70���Ƿ�_ZER �*��s��G� @"���~�O/ RI���
����ɠ�����'�L����T`�W ATUS�p�C_T����O�B+pY�B���3�.�0��� D�e�N� LҾ��M��!��o��XES���һ҆���1�����R�UP:��0��1PX�y�b��3�ǂ���PG텳>��$SUBA�~���AA��JMPWA�IT��r�Y�LOWp/�^�' CVF��vc�\�R���q�C�C��R��i��IG�NR_PL�DB�TBW P�1d�BW� ���U*��IG�L��Ic�TNLND����R֡5B�PN��E�PEED��T�HADOWW b����ES�M�b�+�P0SP]D��� L��Ar�0Q0m�/�{�UN �dy���R�м�LY0���K�_J2�P�H_PK����RETRIE��i��'����FI��� �:����� 2}���DBGLV��?LOGSIZ��1KKTy�U�s2D8�n �_TX�EM�`!Cn�F�X ARR.R>+�CHECK��1���P��p�c������LE�4pPAB#@T��C�O��P��p�bAR%"�Ј�#�1'�O� 0��`ATT���x�%X ��1��UX���sPL,  $��~/QSWITCHT�Z�aW�AS����SLLBp��_ $BAv�D
C2�BAM�����э�J5L���6|�|_KNOW�4���U=�AD��`�x�D��)PAYL#OA��@%#_��.'T�.'Z+#L�AA�qމ0LCL_ʐ !�pg"�Ӂt$˲�&F�)Cgpb*�e$�`Ib(Ripb'{��~$B7`ʑJE��!_�Jl!��֑AND�z�U�
4l"�!(�"aP�L�AL_ �@`x�ѐ����PC>�uD*#E=��J30�36� T�`PDC�K�22�CO�p_�ALPHC3�3BE0БsaC?U<2��b��>� � �.�$/WD_1+*2U$D�pAR��H�5FC塯TIA41I51I6>�MOM��=C]CJCh]CWC�Bp�AD=Cp�FJC�FWCPUB�RbD�EJC�EWB'�@�30ʑq�  �� MO"L� ��*�T���� e$PI����3���0'&Y��J)&YI2[I@[INS�DS�V�V�ޠ2������1�HIGo1�q�j��V j�q�����V�S�X��x�Y��q�SAMP�Ѐ��:d�W;cq�3 Q�iaʐS�Œxd ��fj��0�i@Œߠ �:@�e/0��H��cIN�l/0c�h�k�d�q��jx�d{2{GA�MM�eSU�A�$GGET�R��3�D�4v҂
$60IBR�Ѻ�IL�$HI:�_�����Œ�vEѐ�xA�~�p�vLW�}�v�|��y��v�2�V�51C���CHKİ��q�x>I_`�ޔ.2�8 .1�e|�uCޔ�F{�33� �$e8 �1��I�RCHk_D����RNs�8���LE���R�����8Ѐ��MSWF�L���ASCR�1#00{�. xd39]���gʐ=@�iq�j���P�I3AVMETHaO�æ��妒AX$����X4�p�ER)I��:d3fsR�� 5�	�Q�0FWt;ac$��c�(�L�;a=�OOPa֑S��aN֑APP��F�`� W�x�c��cRT��2�O0j�0�������DR 1�%��D��ѪlNPѢRA� MG���TSV	Q��P; CURC��G�RO7���S_SA��ܴ5���NO�0C �����45��t�?6/H/ TX����zP��UϸCDOi�A�rdyes� �e�X��W��X3�/Ŭ�k# �DMU�o � ��YL$S�!�g��S�"6A9��K���!�����!�_�C���M_W�d���C�����?�M@���ˇ ��21~�L��T�K�� PM&�R�C �}�R��WE�S$��L3X!E� �4Cү4CҶ4C�W4����pN��sf��/0X��O�3.1Z�� P{�T� ���M�� z�w���������4@������ �� P�1_Z� |v1��5�]I��JC ��WC5�6J���PJu�uM�s��� ��@q�P��PMO�N_QU?` �{ 8� QCOU��nQTH_�HO~�n:�HYSES�F:�UE%�+��OX�  ��P#ПuV��RUN_TO��q g�R
P� P! ��C����IND}E�ROGRA���J��2C�NE_NO���IT�A��g��INFO��� �b������ ��I���� (SLE�Q�V"�U" ����S�U��� 4� E�NABqҁ�PTI�ON
�ERVE��R~�Q�VGCF._� @.�J �.1V����pR�x��B�@EDIT��'� �R���K�A�S5�qE�pNU�AUTQ�	COPAY�A�P*�Q]�M�q�N48M�PRUT�R ;N� OUC��Q$G����R�GADJ��� hv0X_��I���п�пW�P�����S��rN0_CY�Cq��RGNSr[�s�=�LGOZ���PNYQ_FRE�Q�BW�`�VP!SIZn[�LAœG!�8XC�`�UCRE�p��f[�IF@Q��NACa�%�$_GœST�ATUv�œy�MA�ILAb�1�!
�5�L�AST�!�1"$EL;EM_� �\�iFEASIl3�nb g�Z�2��>�96���`�pI����G"�Q=� �L�n2ABU�0E��r�PV�!�6BAS�2��5�r�AU�P�PJ��$�1�7RM�@R h3Ł���3���P�r�!��4Q$"S�~�	~E2 2� �c ���d+F�2*G�2"Э`���2VGW�DOU�����r�"$P �@Ҟ)GRID��U�B�ARS�WTYm ��д`O����� �t�_�$!��B�DO|��\� � ����POR���C���C�SRV� )TVDIS�T_�P4PFT�P�PW�PPW4NY5NY6JNY7NY82Q�Fbr�_�r�$VALAU�3(�+4)0�F[�� !hL���b�C�!%���AN'���R�!��T")1TOT�AL_�$l06bPW�=#I�AKdREGENIj^b��X�8��=�� f �TR�3�"IaC_S+��g^`��V���b��2E�# �?�p(2�� cV_H�@�DA ��`pS_YhY���a&S8�AR ��2� �IG_CSE6�`R�%_��v�dC_�F$CMm�,f�wrDEh�?p�r�I]�ZvsPsq!�RE�NHANC&�� pAj�"d#qGINT1P��F}���MASK퓸0OVR��� �<�!Ł �Gy�R��D�d�O�J6�k�F�PSLG|Hp�Q� \ 1� b%Z�$�3`� S���$�qUY�y����cd��ZQU�Aw�TE��>@� (�a�JV�Q�q#IL_M�p$�Vt2����TQ� ����0C���VB�CP�P_�J�Z�mMq�V1p�V1~�U2��2~�3��3~�4��4~�� ��<������IN�VIAB0�J�7��>�2:�U2F�3:�3F�4:�4F���Y�r�U��gP�
�tP��'��PL�� TOR$��IN���u�5����T $MC_FC�X��LC�B��u�)`M��I�s*�rC ���)�r��KEEP_HNADD#��!e��0o�C�ѳ� ���A$�����O�d��>"��`���w��REM�����!�Bµٱ�޸U�$e��HPW�D  e�SB�M�q�@COLLAAB"��P��'a�" cIT' ��INO)�FCALh�
���ܛ ,��FLnб1O$SYN���M���Ccr��`UP_D�LY���r�DEL�A���!�"Y �AD� �.�QSKIPNG�� �
P��O��˂K���P_����� ������#��#� gP"�tP"ځP"ڎP"�ЛP"ڨP"�9��JS2R ���dX�0TJ#����)1�Ѭa�p����a�R RDCa.w�� �� R���R�!�=��-DRG�E� W3�{BFLG��0��SW{	-DSsPC��!UM_�о��2TH2NuA���� 1� ������A[ �� D���x]�02_PC���S���1Q L10_Co"����q ���JPٰ 7��6K�+��� �.�NE���N���b\r�3RC���p��}��DESIG��.JEVL1��1��k�v��10ٰ_DS��K�j��`C11��� lV�������iI�AT����AS'J N$	C�
���oHOME4 ��
��2������� P2D����3���g�y���� 
��4�����L,> ����5���as����V6�����//&/�8/ K��7����[/m//�/�/�/ x��8����/�/�/X? ?2? ��S)�>���  �1���s`Y�V۰E�D�� T���4,f�3IO���
II�0XrOe�_�OPE.C&b�3�P�OWE�� ��0������&d ��}�eB$DSB���GNAr�%c��Cx���Q�S232�5'� ��Z5��׀�ICEUS/cSP�E���QPARIT�q$aOPBQ��RF7LOWApTR�01b�UJsCU�@6��Q�UXT�q�Q�pER�FAC�DʰU `�VSCH�Q� �tV��_�@kpc��$�`�`OM*p��Ap>�#�p%�UPD<�����aPT�0|uEXhЙX|S!%�FA?���r��q�a � ����`;b K�AL"$� ��U��]B�a�  2� �S����0�	� �$t{�����GRO�`�*dT�(p6fDSPBfJOG�`�C����AZ�N������z"VK�P_MIR^a�~d�MT3��cAP@%����`}t��Sp��`R��
��eBRKqHUQ�V��AXI�1  �bc�r-b�qx9�7e�`BSOC6f�۰N2uDUMMY{16O�$SV���DE3A�CF�wK�20�D�pcOR{ws0�N�p|vFp�w[`O�V^eSF�zRUNĴs�rF�vQ�cUF�RA�zTOTLC1H�����OVlt[�[`WP�7�[c���r?pr��_�p� @h�TINVEG@n1O�FS\�C�P�WD��q��q>qf2�eXpT�Rr��1a�E_FyD�aMB_CW�
��B��B�*��ałˁ?�epV9Q��P&�d�írGƇ�hAM�c`��VP�F�!�_M݀0R_�CS�T$���|�Q�3T$HBK�Q,�fm�IO�5|�&A��PPAp��������,�&BS�DVC_DBъ0ސ�Q�Bސ�7�Q������F���3���L�E���+P�`lqU8�3P`FCAB�Ё2@~㷀8û` ���O��UX�fSUBCP �[�-��/��P�/Ѯ�ރ�bB��$HW_C��	P/ы���?�q0#��P�$�UP�t	��AT�TRIh��h`CY�C��g�CAB��cF�LTR_2_FI��3�IH��F��PtkC{HK�_SCT�cF_�F_�����FS�A��CHA��}�ֱ�RղRS�D���Aq�S�A&@_�T�}�.���PEM�0��MsTò/��P�ò��K�DIAG~�URAILAC���M`LO"p��Hv�_�$PSNb�2 X��L��PRߐS}�JI���Cёf�	E��FUN��*QRIN1�}�|0^���Q�S_;`��X����0pf���P�f�CBL�Є�.�A'�#�*�#�D�Ap��h�.�'�LD@yP`p����Ca������TI�°���P$CE_RIAa�V�BAF��P�A��,~���T2}�C�S��؁OI����DF_aL�0�r�Q�PLM�}F^�HRDYO�af�RG��H���a|0|p�/�MULSE�p����Qp�$Jxz�J�r�w�{FAN_�ALMp���WRN��HARD�0�VZ0	P]R�2���A��eY_��fAU�Rȴ~RTO_SBR&E��O`#��ӓ��;�M/PINFQ��N�܆�Y�REG�6NV��Pf3�fDA@N��F9L����$M�Ѕ��`S����P����C�MѐNF-��1�h��h��A��0$�1g$Y oQb|�Q�0�� ��c�EG�0+c`p+AR=`CHu25Rr:T���eAXEEgROBnBjREDBfWR,�2 q_�$sSY�`etp�S�WRI,�>�STr@CcPpJ�pE��0G6RrD��;`B� R��7��.2�OTOi��0��ARYBc4~�2�<"�t`FI�`�c$LwINK�GTHSM�PT_�R�F98Rr|XYZ�R��9�OFFZ�S�{o8B@`��`�/�P�P�FI1������CXt��Zd_J�A�R�r`����30Rr�@�*!m�2b"CFA�eDUn�Hu�3����TUR��X�ӛ%BI�X� `�J'FL|�a�8 � ���	3ʡg� 1��0Kg`M�d�&Qs������°�pSORQ@&�Oa�P(���`O� ��1ɐj4��Ma��~4OVE�1MIPk1�� �5�5�6_Q�7c��7��4ANڡV�1 ���1�`�0�k1�5��1�7(E(E�3OaE)Rla�	��E,��P$��fDAA�P���`!�@o�l�o�AX/� �Ro�2��U�EQ��I {��I���JN �J�J@$�J��J��J1[  �F/��I/��I/��I/� �I/�Y/�Y/�(Y/��8Y/�HYeQYYDEBUڣ$����I�	ao�wABo�m��q39Vb�٢ 
$b� LeʡXgQqXg��Xg NXgXg$Xg�Xg����g ��U�LA�B�J5֠�GR�O[�J"��K�B_ /�MF��s� �v5qpK51u�=vAND0���[DL��^A�zw  K���� �x1ѝxN��NT��#��pVEL�5��4�qm��x9��NmA��V�$���ASS  �����* *  ��_�SI@��]#��)�IY�xn��(�AAVM���K 2 T�� 0  G�5�������.�� ��	݀΍�* U��ߏ��!�͌@�L�܁R�����̡�e�BS�1  1�6�� <u����
��.�@� R�d�v���������Я �����*�<�N�`� r���������̿޿� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߎߠ߀���������߱��pM�AX/� ���nʓ  d�IN��*��PRE_EX�E;�g�J�!43��|T�e�IOCNV�"<� �&�P��a ;��Ɨ��IO_�� 1]r�P $b���0��V���U�?���� �$�6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o(:L^p ������� � �$�6�H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z��������ԟ����LAR�MRECOV �~�!�J���LMD/G ���� ��LM_IF  ��+��ߥ���ɯۯ������0�B�S�, 
 S�|���� ����ƿؿ�$��� ��1��U�g�yϋϝ���NGTOL  �~� 	 A �  �����PPI�NFO Z�� Y��*�<�N�!�  f�P�~�?�mߧ� ���ߵ������%��5�[����χ��� ����������)�;��M�_�m�PPLIC�ATION ?����H��HandlingTool ��� 
V9.10�P/30��j�
�88340����Fy0����1028���������7DF1x��j���Nonej��FRAj� �6w�_ACT7IVE�  �����  �UTOM�OD� ^��ÊCHGAPONL�� �OUPLE�D 1��� �
 2�CUR�EQ 1	��  UT<<<	����@��<����H�k�HTTHKY�A�o��� ////�/S/e/w/�/ �/�/�/�/�/�/?? +?�?O?a?s?�?�?�? �?�?�?�?OO'O�O KO]OoO�O�O�O�O�O �O�O�O_#_}_G_Y_ k_�_�_�_�_�_�_�_ �_ooyoCoUogo�o �o�o�o�o�o�o�o	 u?Qc��� �������q� ;�M�_�}��������� ˏݏ���m�7�I� [�y��������ǟٟ ����i�3�E�W�u� {�������ïկ��� �e�/�A�S�q�w���NTO����DO?_CLEAN����NM  �� <_�qσϕϧ��BDSPDRYRLϊHI� ;�@L� �%�7�I�[�m�ߑ���ߵ������߇MA�X~�������	�X����PLU�GG� ���PRUC��B9�=�����c�Oh�����SEGF� K������9� K��%�7�I�[�����LAP�������� ������	-?Q�cu��TOTA�L+�T��USENU��� ޸���NRGDISPM+MC��0�C���@@���O�������_STRIN�G 1
�
��M� S�

~^_ITEM1h  n����� ���//&/8/J/ \/n/�/�/�/�/�/�/�I/O SI�GNALbT�ryout Mo{deiInp0�Simulate�dmOut,<�OVERR�� �= 100lI?n cycl 5m�Prog Ab�or63m4St�atusk	Heartbeatg�MH Faul<�7�3Aler�9�/ �?�?�?O#O5OGOYOkO}O ��d�� v�O�O�O�O__(_ :_L_^_p_�_�_�_�_��_�_�_ oo�OWOR��dJa�O$oro�o �o�o�o�o�o�o &8J\n�����~POb�1�p bk��#�5�G�Y�k� }�������ŏ׏������1�C�U�g��rDEV�~������˟ ݟ���%�7�I�[� m��������ǯٯ�|���PALT�M 6�bo�^�p������� ��ʿܿ� ��$�6πH�Z�l�~ϐϢ�$�GRI�d��N���� �&�8�J�\�n߀ߒ� �߶����������"�4�F���� R�M~��� X��������� �� $�6�H�Z�l�~�������������l�PREG:�# ����J\n �������� "4FXj|�~�-�$ARG_J`�D ?	������ � 	$�&	[�]���')��SBN_CONF�IG� �$1#2�=!!CII_SAVE  �$F!9#��TCELLSE�TUP �%�  OME_IO��-�,%MOV_qH� �/�/REP����/�UTOBAC�Kv!�@"F�RA:\ X�/F '`�0�C8� T;?  �23/07�/18 17:5/0:04(`�?�?�?�?4<��O�6OHOZOlO~O�O� $O�O�O�O�O__�O <_N_`_r_�_�_�_3_ �_�_�_oo&o�_Jo�\ono�o�o�o�o����  /1_3_\A�TBCKCTL.TM���o+=.;INI9�v56%�J!0MESSAG�V dqF!�o{ODE�_D� Y&6%�xOx���3PAUS�� !�� ,,		� ��� �4��@�B�T���x� �������ҏ�����B����t�pTSK�  �}C?I0UgPDT�pbwd����vXWZD_ENqBbt2*��STAau�����XIS$ U�NT 2�C!�E � 	 m��oRo����(��� r��ߧ�
�����Y!k89�r����F�Бv�+��3�p 0 [?]= 8�a�¯p��������MET��2i�b# P�A�ϴ�Am�xA�R�7;_@���A�?�٭�>a5o>ٹ��>p��5�%�>B�
>H����SCRDCFG� 1�%1 �^%C"篻�Ϳ@߿���<?
QZ) ��e�wωϛϭϿ�&� ��J���+�=�O�a�0��߼1GR���X����`NA� �s	4��_ED`p�1��� 
 ��%-�`EDT- ���*�B�]�b?$� Q-3�
"Ox�&
��  ����!2��#� �G�f5b���G����6����3 ��+]���̔\�� Z�l�����4K�� �����t�&8�\��5�d����@���(��6 �S0/w��/w/��f/���7�//�/ C/���/C?�/�/2?�/B��8{?���?�f����?OV?h?�?�?��9GO�?�O�?i��pO�O`"O4O�OXO��CR�� �/__q_ =:_�_�O�O�_"_����NO_D�EL�ߞ�GE_U�NUSE�ߜ�IG�ALLOW 1���   (�*SYSTEM*�֣	$SERV�_GR�k_`�pRE�Ghe$�c֬_`N�UM�j�c�mPM�U`֥LAY��֬PMP�ALap�eCYC1�0�^�n�`�n%sULSU�o�mr�qjc�L;ttBOXO{RI�eCUR_ap~�mPMCNV�f�ap10~�pT�4DLIǐZ|i	*PROGRAgdPG_MI�n��)�AL�u6� ��)�BT�_n$FLUI_RESUw0���o��ÄMRvn�`�\�_Β��+�=� O�a�s���������͟ ߟ���'�9�K�]� o���������ɯۯ�����#��RLAL_?OUT Nk�����WD_ABOR�p/o��ITR_R_TN  �D���~��NONSTO����� 8hCE_R�IA_I,`��������FCFG� ���ĨN�_�LIMvb2��� �  � 	���gϳB<�҄��e��@� VϷ�����¨H
��ߒ�2�PA�n�GP 1�ޥ�n߀ߒ�QܟC>  C.���f���z���߶Ї�Б��Ж�Р�Ъ�д��Թ�����������C}���ǀ CѶе�J��G?��H=E�PONFIπ��nd�G_P�p1;� �U;ծ������������,�d�KP7AUS~q1;��� �r.�t�;�b��� ������������0 @fL�����6�M��NFO 1�?�� ��T��B�̵���5Au��9	�]�Ǝ��@��K D�5Oy���C����($6�T5+��P�� 8�h��Ca��.~:���1５��O�ϨG���COLLECT_��?�x�ǯEN��p������NDE��?�;c�R�1234567890'�Bya�//&��HC��C)j/�/y\ i/{/�/z[�/�/?�/ �/?`?+?=?O?�?s? �?�?�?�?�?�?8OO O'O�OKO]OoO�O�O@�O�O_�O�9��� ��IO #!)������_��_�_�_`WTR6�2%"D](�{Y
�O�^�o�#o] jt�i_�MOR9�$;� �|�B��.`�e  �i�o�o�o�o�o�kbbT1�:�%pm,t�?]�]���>q�KFt�
`�R�&�utqtr�C4  A���Ț�x�A����BʤpCd B��d C7  @�r��q�:d�QbZqI#'d}?�s9�(pm����}dZqT_DEFB� {%oR��thPNUSE��s���g��KEY_TBL � ������	
��� !"#�$%&'()*+�,-./(':;<=>?@ABC)��GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������,��������������������������������������������������������������4Q��L�CKp�ٹ��p�ST�A���t_AUTO�_DOζkv�I�ND�ٞ�R_T1���T23�ݵʳ���TRL(�LE�TE��z�_SCREEN ;ڿkcsc�U�ʰMMENU 1)l� <7�@�� ����F��#�I��� Y�k��������ſ׿ ��6���l�C�UϢ� yϋϱ������� ��� 	�V�-�?�eߞ�u߇� �߽߫�
������R� )�;��_�q���� �������<��%�r� I�[������������� ��&��5nEW �{�����" �X/A�ew�����/)\ʠ_?MANUALo�*��DB'a.b����DB�G_ERRL.�9*֫�Q /�/��/�.L!NUMLKIM���lu
L!�PXWORK 1+֫�/#?5?G?Y?|k?mDBTB_��G ,{-�s�Qst�3QDB_AWA�YT#�QGCP �lr=���"�2_A!L� ٟ�2P"Yn���tlpE(_n  1-�[,p
?POJf@O}O6�6_M�IS֐�;�@�p�CONTIM6���lt��FI�
� CMOTNE�NDt�DRECO�RD 13֫ y��OxsG�O�KQ 9_x{�2w_�_�_�_DX �_�_K_ oo_$o6oHo �_�_~o�_�oo�o�o �o�o�o �oD�oh z���1�U 
��.�@��d���� �����Џ�Q��u� ���N�`�r���󏨟 ���;����&��� J�5�C������ȯ 7��ׯm�"���F�X� j��y����Ŀ3�� ��ϣ���Bϱ�f�տ �ϜϮ���[���S�߀w�,�>�P�b��Ͽ2TOLERENC�4sB�B�0L��L �CSS_CNST_CY 249�Y 	e�B��������� �#�5�G�]�k�}�� ����������������DEVICE ;25�� �6o� ���������������&�O��HNDG�D 6�۬0Cz�9
Q��LS 27Y�8������:��PARAM 8,I�2�5&��ySLAVE �9YE_CFG� :F&d�MC:\��L%0?4d.CSV%@�c�B�A �C	H kkO&/B/
X�&2"_!o/])<\!1@JPя#N.�A�1n_CRC_OUT ;Y���1*_NOCOD�z<,G�SGN� ="UR#M��18-JU�L-23 23:�46�0A:917:�51�~� V�hr9n1&o061��M��Þ�ǧj��1�>�VE�RSION �):V4.2.�11�KEFLOG�IC 1>�� 	�(1@I�!M��2PROG_ENqB Xa=CULS�G� `�2_ACC�LIM�F����|CWRSTJ�NT�G
S���1MO�FLX!2�DINIT� ?��"U�� �FOPTu ?	��F�B
 	Rg575&'P74,Y56-X7-W50QX�4�WR2-T�({_�7
TTO  ]�?�_�6]V�@DEX�Gd�B�� �SPATH ;A):A\�_5o�Go|�HCP_CL?NTID ?�6� �+Ӈo���IAG_GRP {2D� �� 	 D� � D�� D � B��Т��f�f�j�`���o�l�a����%��B��N�C�-BzBp��e`��imp2m7� 7890123�456xq�G�`� � Ao�
A�j{Ad�]���AW�AP���AJ=qAC3w3A<�4z�jL�p�!@��]pA�q���A�����B�4�lf�dX�!
��ru�ppQ�Aj��HAeG�A_��pY��AS�pM�2�F�RA@(� �J���t�J��I��@�p��������@��HL�^�p���������33<���=q@~�R@x�Q�@q�@k��@dz�@]��Vff؏����� ���s>�l��@�e@^J�W
�=@Pv�G�@u@v�7ڐ.{d��v���������S>�M����AR�<(�@�5Ґ/\)@(��@!R�֏ �� $�6��ĭ���ܯ"� 4����V�|�Z����� <�N�������0�B� ̿R��B�`�r5���M�xّe��m>��R���?�33?9���{���m7'Ŭ���6��4�F���L�m@ž�����ڐ␀N�Њ=@V�pAh�����c�= c<��]�>*�H>V�>�3�>���~�m<���<b��a�i�L. �?�� �C�  <(��UX" 4� >��ё��ٝiA吳 ?�el���t����,� �H��8�b���r��z�x����x�?�7���>�(�>!�����=����m��G��G��m�����I��m����i�@��Ҁ�@Q�?L ��Ly�o�g�v\����]p'�@����8����	�gC� �̇�Cu��Zl �<� ���`��&%�18� �����4J�6�<�D5�OL��rC��� >T&U�Q���$�z�	��($6�T��Á�i���x�������=ʝm;��t���9/�aCT_CON?FIG E?i3�eg�%�aSTBF_TTS�G�
UI�#�0�C�A�&�� MAU�@JOJ"M_SW_CFX F�k�  �p�:OCVI�EW� G�-�a���o=?O?a?s?�?�? �B+?�?�?�?�?OO �?>OPObOtO�O�O'O �O�O�O�O__(_�O L_^_p_�_�_�_5_�_ �_�_ oo$o�_HoZo lo~o�o�o�oCo�o�o �o 2�oVhz0���@,RC�#{��"!L�~���A��0�e�T����$SBL�_FAULT �I�z 8��GPMS�K�'��L TDIAOG J\)�!���1�UD1�: 6789012345�p"1�j'�uP&/O�a�s����� ����͟ߟ���'� 9�K�]�o�����y���
>���F&TREC	P���
���%��� =�:�L�^�p������� ��ʿܿ� ��$�6πH�Zρ�������7U�MP_OPTIO1N� ����TR�"�#:����PME�%���Y_TEMP  È�3BȞ �1��A.��UNI�� �%1��&YN_B�RK K?6EDITOR����
���_ԠENT 1�L�y  ,&�PART1 T�LOG ���߫�&MAI���߫����2��0�&�OMAY�[�  D��߇�n�� u����J���n�
IRVW�AI����&-BCKEDT- ���/�f�PICKSIM_��[�f�y���o"�x��������� ����3WiP �t�������~�MGDI_S�TAD� !1�y�NCv71M�+ �`�(r��
��d��� ��/!/3/E/W/i/ {/�/�/�/�/�/�/�/ ??/?A?S?��j?|? �?�?�9��?�?�?�? 
OO.O@OROdOvO�O �O�O�O�O�O�O__ *_<_�:c?m__�_�_ �?�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/A[_ ew���_��� ���+�=�O�a�s� ��������͏ߏ�� �'�9�SA�o����� ���ɟ۟����#� 5�G�Y�k�}������� ůׯ�����1�K� ]�g�y���A�����ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�C�U�_�q߃� �߯����������� %�7�I�[�m���� �����������!�3� M�W�i�{����߱��� ������/AS ew������ �+E�Oas ��������/ /'/9/K/]/o/�/�/ �/�/�/�/�/�/?#? =/?Y?k?}?���? �?�?�?�?OO1OCO UOgOyO�O�O�O�O�O �O�O	__5?G?Q_c_ u_�_�?�_�_�_�_�_ oo)o;oMo_oqo�o �o�o�o�o�o�o �_?_I[m�_� ������!�3� E�W�i�{�������Ï Տ�����7A�S� e�w��������џ� ����+�=�O�a�s� ��������ͯ߯�� �/��K�]�o���� ����ɿۿ����#� 5�G�Y�k�}Ϗϡϳ� ���������'�9�C� U�g�ߓ��߯����� ����	��-�?�Q�c� u����������� ��1�;�M�_�q��� ������������ %7I[m�� �����)�3 EWi������ ���////A/S/ e/w/�/�/�/�/�/�/ �/?!+?=?O?a?{ m?�?�?�?�?�?�?O O'O9OKO]OoO�O�O �O�O�O�O�O�O?_ 5_G_Y_s?�?�_�_�_ �_�_�_�_oo1oCo Uogoyo�o�o�o�o�o �o�o_#_-?Qc }_������� ��)�;�M�_�q��� ������ˏݏ�i %�7�I�[�u����� ��ǟٟ����!�3� E�W�i�{�������ï կ�����/�A�S� m�w���������ѿ� ����+�=�O�a�s� �ϗϩϻ�������� ��'�9�K�e�[߁ߓ� �߷����������#� 5�G�Y�k�}���� ���������1�C� ��o�y����������� ����	-?Qc u�������� �);Mg�q� ������// %/7/I/[/m//�/�/ �/�/�/�/?!?3? E?_i?{?�?�?�?�? �?�?�?OO/OAOSO eOwO�O�O�O�O�O�O �/__+_=_W?I_s_ �_�_�_�_�_�_�_o o'o9oKo]ooo�o�o �o�o�o�o�O�o# 5O_a_k}��� ������1�C� U�g�y���������ӏ �o�o	��-�?�Yc� u���������ϟ�� ��)�;�M�_�q��� ������˯E����� %�7�Q�[�m������ ��ǿٿ����!�3� E�W�i�{ύϟϱ��� �������/�I�S� e�w߉ߛ߭߿����� ����+�=�O�a�s� ������������ �'�A�7�]�o����� ������������# 5GYk}������� �$ENE�TMODE 1N�B�� + �������� RROR_P�ROG %�
%���an<TABL/E  �L�����<SEV_�NUM 
  �� <_�AUTO_ENB�  (9_N�O! O�� "  *�Y �JY �Y �Y  +X �r/�/�/2$FLTR/0&HIS����++_ALM 1P.� ���Y,��+�/2?D?V?h?z?�?�/_�8   ��W!�:� TC�P_VER !��
!Y�?$EXTLOG_REQ�&s�))#CSIZ,O�DSTKIIG%�� BTOL  ���Dz�"�A D_BWD�0�@�&زA#�CDI�A QB��C���KSTEP�O�O� >�@OP_DOkO��FACTORY_�TUN�'d3YDR_GRP 1R�	�!d 	�?�_{P��*u����RHB ��2� ��� �e9 ����V{S�_�]�{PB���B���]C��B����AԂ=B�X���]A��B�^�B�]gA����AI��B�V�]�_WoBo{ofo�o�o�o�o  @��:A|=@9�q��o��
 Fǂ5W&b�`��A�>��o	2�o�o\G܀�]�  �qA���`�33�r�33^�]@UUT�z@�`��pj$>u.�>*��<����]�E�� F@ ��p&��]J��N�Jk�I'PK�Hu��IP�s�F!���]?� � j��9�<9��896�C'6<,5����~���=����a��� �_&����#tFEATUROE SB��@"�Handl�ingTool �	���Engl�ish Dict�ionary�4�D St��ard�	��Analog� I/O@�I�gle Shift\��uto Soft�ware Upd�ate��mati�c Backup����ground� Edit��C_ameraW�F[��CnrRndIm����ommon �calib UI���n͑�Monoitor&�tr�?Reliabp���DHCP�]�at�a Acquis�5�^�iagnos���T�x�ocume�nt Viewe�A�`�ual Ch�eck Safe�ty!��hanc�ed!����sʠF�rސ�xt. D7IO 1�fi��&�wend��Err@�QL��B��sA�rR��1� �@�FCTN_ Menu�v\����TP In��f�ac���GigE���εƐp Mas_k Exc��g#��HT��Proxy� Svˤ�igh�-Spe��Ski��Ŧ�5�mmun�ic��ons<�u�r����s�X���connect 2s��ncr��struH#�qʚ�e��۠J����KAREL C�md. L �ua����Run-Ti�"�Env�Ȅ�el� +��s��S/W��License�ݣʬX�Book(System)�MACROs,3�?/Offsew�V�aH5���q�[�MR:��6���MechSt�op�t����V�iS�s���x��T������odq�witch��ߚӡ�.{��Op�tm,���fil�ʬ��gi�V�ult�i-T��Г�PC�M fun�Ǣ�o���ޢ����Regi�K�rW���riàF�����U�Num S�el��� � Ad�juG��=�s�N�t�atu��f�Ū�R�DM Robot> �scove)����ea��"�Freq� AnlyW�Re�m��5�n7�����S�ervo5���S�NPX b�x�SN��Cli¡%t��Libr(�E�� ���W o0�t��sGsag����0 ���n���0/I���M�ILIB��P OFirm���P���AccǐϛTPT9Xm��elnn����jղorqu>q�imula?��bu�PaѱƐtZ�(�&�ev.�抐ri۠:USB port ��iPL�aà�R �EVNT��nexcept������X���VC�rR�I���V��o"�%W�z+S8 SC4�/S�GE�/�%UI�Web Pl}� >�i�'4�����x�ZD?T ApplP��x&?|7Grid��playv=� ���7Rf".7��6���/Y��-10iA/8L��?Alarm �Cause/��e}d*�Ascii��<�Loadʠ:JU�plP@�l�7�G�u=�rO�BP��Ֆy�cp�����蠕�R�A� �9�NRT�J�On�e Hel��漿��������1tr;�ROS WEth
�t�BeW7�iR�$2D Pk,;�uVIm+�Fd�� ��^nsp���Q�6�4MB DRAM��O�SFRO�_ېe3llW��shao" gcK�e��p�2ltyp�s'�ԗ�B��:D�.�maiܠ;P�T�qV�R7�:�FL!PSup�c�p�� pL���cro~����W�4��&��auestz&rtڡ���/�3DL}|�Q����Ty,K��l Bu�i��n�/APLCd��uVZ��/CGl�N�CRG#��$D���@�R�LS[��%BU�w��%Kі��!TA����B�,يE�TCB��ʏ��/��^�TC��v��%��TEHǟٖ"�BؗV�����/��F�H����G:���n���d����H¯��IA߯��ޯ��LN���M@��D���D�����N�B��P��������RR�B��Sڿ�����W.�8@Ǣ��$VGFf�x�P2Z���2��ǂϔ�IB�ϔ�D�ϔ�Fr������"TUT��0�1J�\�2f�\�TB�GG��rain��UI*ЦUHMI��r ponU2�8��af{ �R�v�VKAgREL��_TP� �e��R9�0�B�o� f�x���������� ���5�,�>�k�b�t� �������������� 1(:g^p�� ����� -$ 6cZl���� ����)/ /2/_/ V/h/�/�/�/�/�/�/ �/�/%??.?[?R?d? �?�?�?�?�?�?�?�? !OO*OWONO`O�O�O �O�O�O�O�O�O__ &_S_J_\_�_�_�_�_ �_�_�_�_oo"oOo FoXo�o|o�o�o�o�o �o�oKBT �x������ ���G�>�P�}�t� ������׏Ώ���� �C�:�L�y�p����� ��ӟʟܟ	� ��?� 6�H�u�l�~�����ϯ Ưد����;�2�D� q�h�z�����˿¿Կ ���
�7�.�@�m�d� vψϚ��Ͼ������� �3�*�<�i�`�r߄� ���ߺ��������/� &�8�e�\�n���� ����������+�"�4� a�X�j�|��������� ������'0]T fx������ �#,YPbt �������/ /(/U/L/^/p/�/�/ �/�/�/�/�/??$? Q?H?Z?l?~?�?�?�? �?�?�?OO OMODO VOhOzO�O�O�O�O�O �O_
__I_@_R_d_ v_�_�_�_�_�_�_o ooEo<oNo`oro�o �o�o�o�o�o A8J\n��� ������=�4� F�X�j�������͏ď ֏����9�0�B�T� f�������ɟ��ҟ�� ���5�,�>�P�b��� ����ů��ί���� 1�(�:�L�^������� ����ʿ��� �-�$� 6�H�Zχ�~ϐϽϴ� ��������)� �2�D� V߃�zߌ߹߰����� ����%��.�@�R�� v����������� !��*�<�N�{�r��� ������������ &8Jwn�������  �H552��2�1R7850�J614AT�UP)545)6�VCAMCR�IdUIF)28neNRE52XwR63SCH�DOCV�CSU�869)04E�IOC�4R6=9XESETAW�J7WR68M�ASKPRXY�}7OCO(3�A! (3`&J6�'53�H�(LC�HH&OPLGA0^x&MHCRI&S�'�MCS@0$'55�4MDSW!7k'OPk'MPRl&��(�0(PCM|R0`g7! 4� �'51L�51�80LPRSv'69`&FRDd�FREQMCN�93(SNBA���'SHLBFM�'G�82(HTC�@TMIL�T{PA�TPTXYF#EL�6� �8�J95�TUTvl'95`&UEV&wUECH&UFRd�VCC XO�&VI�PdFCSC�FCS�G��IWEBn@HTT@R6���HCG_WIGGWI�PGS�VRCdFD�Gk'H7�R66�LR7'R�8R5�3�768�82x&Rڦ*4�W664R6�4NVD&R6��'9 �X�9 �D0:+gF~hCLIP8K�CMS��`@STmY$WTO@NN`&�ORS�&M�8OL��hENDLWS��hFVR�V3D�$X{PBV�FAP�L�APVl&CC�G@CCR�&CD�WCDL�VCSBn�CSK,6CT{GGCTBHV�p�hC(F4�p�xC<WTC|�p�pwTC�wTC&CcTE�9�|wTE��9�0WTF�xF�hGR�xGx�$�H$�IF���$��GCTM�hM��M�xN$�P��P��xR�x�hTS�xW�8��VVGFP�P2F WP2�6e�\�B\��D\�F|VP��VqT��VTB�w-V�IHWGV�P՗K$WV_V��)�;� M�_�q���������˯ ݯ���%�7�I�[� m��������ǿٿ� ���!�3�E�W�i�{� �ϟϱ���������� �/�A�S�e�w߉ߛ� �߿���������+� =�O�a�s����� ��������'�9�K� ]�o������������� ����#5GYk }������� 1CUgy� ������	// -/?/Q/c/u/�/�/�/ �/�/�/�/??)?;? M?_?q?�?�?�?�?�? �?�?OO%O7OIO[O mOO�O�O�O�O�O�O �O_!_3_E_W_i_{_ �_�_�_�_�_�_�_o o/oAoSoeowo�o�o �o�o�o�o�o+ =Oas���� �����'�9�K� ]�o���������ɏۏ��  H�55Ȕ�����R�78�50	�J6;14	�ATU�?��5459�6	�VC�AM	�CRI��U�IF9�28��NR�E�52x�R63��SCH	�DOC�V��CSU�86�99�0H�EIOC�ɛ4(�R69x�EgSETY�w�J7w��R68�MASK^	�PRXY��7	�OCOy�3Y�(����8�3تJ67�53�(�H�LCH��O�PLGY�0��MH�CR��Sw�MCS�X�0��55H�MD�SWٻ�OP�M�PR��(�08�PCM��R07˅�H�l��(�51h�51x��0h�PRSx�69�تFRD��FRE�Q�MCN	�93�8�SNBAٛ�SHLB	�M7��ȼ�28�HTCX�TMsIL�(�TPAH�oTPTXy�EL��ą�(�8'�%��J9�5��TUT�95�تUEVx�UECUFR��VCC�X�O��VIP��C;SC��CSGȚ��I	�WEBX�HT�TX�R6ל��CG���IG��IPGS�	�RC��DG�H�7'�R66h�R7�g�Rv�R53h�6U8h�2��R6�4���66H�R64�NVDx�R6����h�X������D0��FV�CLI�g�CMS�H�� X�STY��T�OX�NNتORSژ�M��OL�EN�D�Lg�S�FV�RH�V3D�짛P�BV��APLH�A�PV�CCGX�C�CRx�CDg�CD�L(�CSB�CS�K�CT��CTB��� �C8�5 ,Cƨ�TC��5 �TCv�TCx�CTE���� �TE�� ��TUF,F�G,G�-
�,H�,I�E0�,��WCTM�Mx,M�UN�,PH<P,R,��TS,W�=(�V�GFKP2X�P2���5@(LB(LD(LF6��VPW;VT��@�(�VTB�V�I�Hw�V5��KK��V ���_1_C_U_g_y_ �_�_�_�_�_�_�_	o o-o?oQocouo�o�o �o�o�o�o�o) ;M_q���� �����%�7�I� [�m��������Ǐُ ����!�3�E�W�i� {�������ß՟��� ��/�A�S�e�w��� ������ѯ����� +�=�O�a�s������� ��Ϳ߿���'�9� K�]�oρϓϥϷ��� �������#�5�G�Y� k�}ߏߡ߳������� ����1�C�U�g�y� ������������	� �-�?�Q�c�u����� ����������) ;M_q���� ���%7I [m����� ��/!/3/E/W/i/ {/�/�/�/�/�/�/�/ ??/?A?S?e?w?�? �?�?�?�?�?�?OO +O=OOOaOsO�O�O�O �O�O�O�O__'_9_ K_]_o_�_�_�_�_�_ �_�_�_o#o5oGoYo ko}o�o�o�o�o�o�o �o1CUgy �������	� �-�?�Q�c�u�����Ы���Ϗ���STD�LANG�� �2�D�V� h�z�������ԟ� ��
��.�@�R�d�v� ��������Я���� �*�<�N�`�r����� ����̿޿���&� 8�J�\�nπϒϤ϶� ���������"�4�F��X�j�|ߎߠ߲�RB=T�OPTN���� �����#�5�G�Y�k�DPN������ ��������%�7�I� [�m������������ ����!3EWi {������� /ASew� ������*� /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?u?�?�?�?�? �?�?�?OO)O;OMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /ASew��� ������+�=� O�a�s���������͏ ߏ���'�9�K�]� o���������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�C�U�g�y����� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� ��������)�;�M� _�q߃ߕߧ߹����� ����%�7�I�[�m� ������������ �!�3�E�W�i�{��� ������������/ASe�h��p����99���$FEAT_A�DD ?	����  	�%7I[m ������� /!/3/E/W/i/{/�/ �/�/�/�/�/�/?? /?A?S?e?w?�?�?�? �?�?�?�?OO+O=O OOaOsO�O�O�O�O�O �O�O__'_9_K_]_ o_�_�_�_�_�_�_�_ �_o#o5oGoYoko}o �o�o�o�o�o�o�o 1CUgy�� �����	��-� ?�Q�c�u��������� Ϗ����)�;�M� _�q���������˟ݟ ���%�7�I�[�m� �������ǯٯ��� �!�3�E�W�i�{��� ����ÿտ����� /�A�S�e�wωϛϭ�����������DE�MO S   �N�D�V� ��zߌ߹߰������� ����I�@�R��v� ������������ �E�<�N�{�r����� ����������
A 8Jwn���� ���=4F sj|����� �//9/0/B/o/f/ x/�/�/�/�/�/�/�/ ?5?,?>?k?b?t?�? �?�?�?�?�?�?O1O (O:OgO^OpO�O�O�O �O�O�O�O _-_$_6_ c_Z_l_�_�_�_�_�_ �_�_�_)o o2o_oVo ho�o�o�o�o�o�o�o �o%.[Rd� �������!� �*�W�N�`������� Ï��̏�����&� S�J�\����������� ȟ����"�O�F� X���|�������įޯ ����K�B�T��� x���������ڿ�� ��G�>�P�}�tφ� �Ϫϼ�������� C�:�L�y�p߂߯ߦ� ������	� ��?�6� H�u�l�~������ ������;�2�D�q� h�z����������� ��
7.@mdv ������� 3*<i`r�� �����///&/ 8/e/\/n/�/�/�/�/ �/�/�/�/+?"?4?a? X?j?�?�?�?�?�?�? �?�?'OO0O]OTOfO �O�O�O�O�O�O�O�O #__,_Y_P_b_�_�_ �_�_�_�_�_�_oo (oUoLo^o�o�o�o�o �o�o�o�o$Q HZ�~���� ���� �M�D�V� ��z�������ݏԏ� �
��I�@�R��v� ������ٟП��� �E�<�N�{�r����� ��կ̯ޯ���A� 8�J�w�n�������ѿ ȿڿ����=�4�F� s�j�|ϖϠ������� ����9�0�B�o�f� xߒߜ����������� �5�,�>�k�b�t�� ������������1� (�:�g�^�p������� �������� -$6 cZl����� ���) 2_V h������� �%//./[/R/d/~/ �/�/�/�/�/�/�/!? ?*?W?N?`?z?�?�? �?�?�?�?�?OO&O SOJO\OvO�O�O�O�O �O�O�O__"_O_F_ X_r_|_�_�_�_�_�_ �_oooKoBoTono xo�o�o�o�o�o�o G>Pjt� �������� C�:�L�f�p������� ӏʏ܏	� ��?�6� H�b�l�������ϟƟ ؟����;�2�D�^� h�������˯¯ԯ� ��
�7�.�@�Z�d��� ����ǿ��п����� 3�*�<�V�`ύτϖ� �Ϻ��������/�&� 8�R�\߉߀ߒ߿߶� ��������+�"�4�N� X��|�������� ����'��0�J�T��� x��������������� #,FP}t� ������ (BLyp��� ����//$/>/ H/u/l/~/�/�/�/�/ �/�/?? ?:?D?q? h?z?�?�?�?�?�?�? O
OO6O@OmOdOvO �O�O�O�O�O�O__>2]  )XH_ Z_l_~_�_�_�_�_�_ �_�_o o2oDoVoho zo�o�o�o�o�o�o�o 
.@Rdv� �������� *�<�N�`�r������� ��̏ޏ����&�8� J�\�n���������ȟ ڟ����"�4�F�X� j�|�������į֯� ����0�B�T�f�x� ��������ҿ���� �,�>�P�b�tφϘ� �ϼ���������(� :�L�^�p߂ߔߦ߸� ������ ��$�6�H� Z�l�~�������� ����� �2�D�V�h� z��������������� 
.@Rdv� ������ *<N`r��� ����//&/8/ J/\/n/�/�/�/�/�/ �/�/�/?"?4?F?X? j?|?�?�?�?�?�?�? �?OO0OBOTOfOxO �O�O�O�O�O�O�O_ _,_>_P_b_t_�_�_ �_�_�_�_�_oo(o :oLo^opo�o�o�o�o �o�o�o $6H Zl~����� ��� �2�D�V�h� z�������ԏ��� 
��.�@�R�d�v��� ������П����� *�<�N�`�r������� ��̯ޯ���&�8� J�\�n���������ȿ ڿ����"�4�F�X� j�|ώϠϲ������������0�  1�6�L�^�p߂ߔ� �߸������� ��$� 6�H�Z�l�~���� ��������� �2�D� V�h�z����������� ����
.@Rd v������� *<N`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/�/?"?4? F?X?j?|?�?�?�?�? �?�?�?OO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �_�_�_�_�_�_�_o o(o:oLo^opo�o�o �o�o�o�o�o $ 6HZl~��� ����� �2�D� V�h�z�������ԏ ���
��.�@�R�d� v���������П��� ��*�<�N�`�r��� ������̯ޯ��� &�8�J�\�n������� ��ȿڿ����"�4� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ߮������� ����,�>�P�b�t� ������������ �(�:�L�^�p����� ���������� $ 6HZl~��� ���� 2D Vhz����� ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ??*?<?N?`?r?�? �?�?�?�?�?�?OO &O8OJO\OnO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_ �_�_�_oo0oBoTo foxo�o�o�o�o�o�o �o,>Pbt �������� �(�:�L�^�p����� ����ʏ܏� ��$� 6�H�Z�l�~������� Ɵ؟���� �2�D� V�h�z�������¯ԯ ���
��.�@�R�d� v���������п��� ��*�<�N�`�rτ� �ϨϺ���������&�5�:�-�P�b� t߆ߘߪ߼������� ��(�:�L�^�p�� ���������� �� $�6�H�Z�l�~����� ���������� 2 DVhz���� ���
.@R dv������ �//*/</N/`/r/ �/�/�/�/�/�/�/? ?&?8?J?\?n?�?�? �?�?�?�?�?�?O"O 4OFOXOjO|O�O�O�O �O�O�O�O__0_B_ T_f_x_�_�_�_�_�_ �_�_oo,o>oPobo to�o�o�o�o�o�o�o (:L^p� ������ �� $�6�H�Z�l�~����� ��Ə؏���� �2� D�V�h�z������� ԟ���
��.�@�R� d�v���������Я� ����*�<�N�`�r� ��������̿޿�� �&�8�J�\�nπϒ� �϶����������"� 4�F�X�j�|ߎߠ߲� ����������0�B� T�f�x�������� ������,�>�P�b� t��������������� (:L^p� ������  $6HZl~�� �����/ /2/ D/V/h/z/�/�/�/�/ �/�/�/
??.?@?R? d?v?�?�?�?�?�?�? �?OO*O<ONO`OrO �O�O�O�O�O�O�O_�_&_8Y�$FEA�T_DEMOIN�  =T�hP��=PPTINDEX�][lQ�PPILE�COMP Tw����QkR�KU�PSETUP2� U�U�R��  N �Q�S_�AP2BCK 1�V�Y  �)�9Xok%�_:o=P �P(oeo;U�_�o o�o Do�o�ozo�o3E �oi�o��.�R �����A��N� w����*���я`��� ���+���O�ޏs��� ���8�͟\�ڟ��� '���K�]�쟁���� ��F�ۯj������5� įY��f������B� ׿�x�Ϝ�1�C�ҿ g����ϝ�,���P��� t���ߪ�?���c�u� ߙ�(߽���^��߂� �)��M���q� �~� ��6���Z������%� ��I�[��������� D���h�����
3�Y��PP�_ 2�P�*.VR:���*�������n �PC���FR6:�4�X�T|P|�y�_PxI���*.FqD/��	�<,�`/�STMk/�/�"�/�-O/�/�H �/?�'?�/�/i?�GIFs?�?�%�?F?8X?�?�JPG�?!O��%O�?�?qO�
JS�{O�O��7C�OOO%�
JavaScrgipt�O�?CS�O�(_�&_�O %C�ascading� Style S�heetsT_��
�ARGNAME.SDT�_��� \�_�U_�A�T�_�_�PDOISP*�_���T�o�_�QNa\oo
T�PEINS.XML�o�_:\�o]o�Q�Custom T?oolbar�oi�PASSWORD�So��FRS:\�#�oD`Passw�ord Configd���<�� ��+�=��a�� ����&���J�ߏn��� ���9�ȏ2�o����� "���ɟX��|��#� ��G�֟k������0� ůT����������C� U��y������>�ӿ b�������-ϼ�Q�� Jχ�ϫ�:�����p� ߔ�)�;���_��σ� �$߹�H���l���� ��7���[�m��ߑ� � ����V���z����� E���i���b���.��� R���������AS ��w�*<�` ���+�O�s ��8��n/ �'/��]/��// z/�/F/�/j/�/?�/ 5?�/Y?k?�/�??�? B?T?�?x?O�?OCO �?gO�?�O�O,O�OPO �O�O�O_�O?_�O�O u__�_(_�_�_^_�_ �_o)o�_Mo�_qo�o o�o6o�oZolo�o %�o[�o� �D�h���3� �W��������@� ���v����/�A�Џ e�􏉟��*���N���r�������$FI�LE_DGBCK� 1V������ <� �)
SUMM?ARY.DG#�ϜOMD:W���ې�Diag Su�mmary����
CONSLOG���p���ۯ���Co�nsole lo�g���	TPACCN�v�%^������TP Acco�untin=����FR6:IPKD?MP.ZIPϿӘ�
� ϧ���Exc?eption$�ջ���MEMCHEC�K��������/�M�emory Da�ta���� l�=)��RIPE��ϸ��'߶�%�� �Packet L<<���L�$�e���STAT!��߯�� %C�St�atus��`�	F�TP�������1�mment T�BD4�`� >I)�ETHERNE�y��f�w�瑱E�thernL�3�figuraCϫ��?DCSVRF(��� �9����� ve�rify all�<���M.c��DIFF1��)���=�S�diff��t�f�>��CHG01�������C����kv�- 	29 2���h�z3���K� �rVT�RNDIAG.LASw(:����O Ope��N� ���nostic����)VDEV�DAT�������Vis�De�vice�+IM�G��./@/�/<��k$Imagw/+�UP ES/�/�FRS:\?\=���Updates� List\?���� FLEXEVEAN��/�/�?���1 UIF EvO��O���,�t)
�PSRBWLD.CMOϜG2#O^?�0�PS_ROBO�WELU���:GI�G�ϾO�?�O��G�igE�(O��N��A�)�AHAD�OW�O�O�Oi_���Shadow C�hange������a�)RRCME�RRa_F_X_�_����PCFG Err{orq tail�_� MA�m�CMSGLIB�_�_�_`so�B6e��|0ico�+a�)_`ZD�O�o\o�o��ZDfPad�o l )RNOTI��o�ow���Notifiqc�� F�AG�� �՟����(���L� �p������5�ʏ܏ k� ���$�6�ŏZ�� ~������C�؟g��� ���2���V�h����� ���¯Q��u�
��� �@�ϯd�󯈿��)� ��M������ϧ�<� N�ݿr�ϖ�%ϣ��� [�����&ߵ�J��� n߀�ߤ�3�����i� �ߍ�"��/�X���|� ���A���e���� ��0���T�f����� ��=�����s���, >��b����'� K����:� Gp��#��Y �}/$/�H/�l/ ~//�/1/�/U/�/�/ �/ ?�/D?V?�/z?	? �?�???�?c?�?
O�? .O�?RO�?_O�OO�O ;O�O�OqO_�O*_<_ �O`_�O�_�_%_�_I_ �_m_�_o�_8o�_\o no�_�o!o�o�oWo�o {o"�oF�oj�o w�/�S��� ��B�T��x���� ��=�ҏa������,����$FILE_�FRSPRT  ��������A�MDO?NLY 1VU��� 
 �)�MD:_VDAEXTP.ZZZ3��䏻�ʛ6%�NO Back �file ���S�6)�����@�	� M�v�����)���Я_� �����*���N�ݯr� �����7�̿[�ٿ� ��&ϵ�J�\�뿀�� �϶�E���i���ߟ� 4���X���eߎ�߲� A�����w���0�B����f��ߊ��E�VI�SBCKs�]����*.VD����U��FR:\��ION?\DATA\��w��U�Vision VD��!�[� m����{��D����� z���3E��i�� �.�R��� �A�Rw� *��`��/� �O/�s/�/@/�/8/ �/\/�/?�/'?�/K? ]?�/�??�?4?F?�?�;�LUI_CON�FIG WU�����; $ �3x�{U�=OOOaOsO0�O�O�I%@|x�?�O �O�O__'\�OJ_\_ n_�_�_)_�_�_�_�_ �_o�_4oFoXojo|o �o%o�o�o�o�o�o �o0BTfx�! �������,� >�P�b�t�������� Ώ������(�:�L� ^�p��������ʟܟ ���$�6�H�Z�l� �������Ưدꯁ� � �2�D�V�h����� ����¿Կ�}�
�� .�@�R�d����ϚϬ� ������y���*�<� N�`��τߖߨߺ��� ��u���&�8�J��� [�������_��� ���"�4�F���j�|� ��������[����� 0B��fx�� ��W��, >�bt���� S��//(/:/� ^/p/�/�/�/=/�/�/ �/ ??$?�/H?Z?l? ~?�?�?9?�?�?�?�? O O�?DOVOhOzO�O �O5O�O�O�O�O
__ �O@_R_d_v_�_�_1_ �_�_�_�_oo�_<o@No`oro�o�o&h�`�x�o�c�$FLU�I_DATA �X����a�)a�dRES�ULT 2Y�e�p �T��/wizard/�guided/s�teps/Expert�o?Qcu ����������Skip G�pance an�d Finish? Setup�D� V�h�z�������ԏ����&h �`.�)`�e!�0 ��2`!��c�aA��ps������� ԟ���
��.�@�R� �2oy���������ӯ ���	��-�?�Q�)e@�)cA�3�E�W�g�rip*pu�ۿ��� �#�5�G�Y�k�}Ϗ� ��`����������� 1�C�U�g�yߋߝ�\� n����ߤ�b�g�%p�TimeUS/DST��?�Q�c�u����������
�?Enable��(� :�L�^�p���������P������ �b�a����������#�24 *������� 1C��y� ������	// -/?/Q/"4F\��$qRegion T/�/�/??+?=?O?�a?s?�?�?�AmericaϿ�?�? �?OO+O=OOOaOsO�O�O�)aym//�O��/�/#sditor �O7_I_[_m__�_�_�_�_�_�_� To�uch Pane�l  S (rec_ommenp)�_ >oPoboto�o�o�o�o�o�o�o�L��O�O5��O	_Racces �?����������,�>���Co�nnect to� Network M���������̏ޏ��@��&�8�J��H�^ !9+=S!_P�Introduct�/�����*�<� N�`�r������Ϻ�̯ ޯ���&�8�J�\�0n������� ��w������YVSafet�A$�6�H�Z�l�~� �Ϣϴ������ϩ��  �2�D�V�h�zߌߞ� ���������߷�ɿ� �[�k�}���� ����������1�C� �g�y����������������	-?[(�5��-�Q� ����"4F Xj|�M���� ��//0/B/T/f/ x/�/�/[m�/� ??,?>?P?b?t?�? �?�?�?�?�?��?O (O:OLO^OpO�O�O�O �O�O�O�O�/_�/3_ �/Z_l_~_�_�_�_�_ �_�_�_o o2oDoU_ hozo�o�o�o�o�o�o �o
.@�Oa#_ �G_������ �*�<�N�`�r����� Uo��̏ޏ����&� 8�J�\�n�����Q�� uן����"�4�F� X�j�|�������į֯ 诧���0�B�T�f� x���������ҿ俣� �ǟ)�;���b�tφ� �Ϫϼ��������� (�:���^�p߂ߔߦ� �������� ��$�6� ��?��c��Oϴ��� ������� �2�D�V� h�z���K߰������� ��
.@Rdv �G��k���� *<N`r�� ������//&/ 8/J/\/n/�/�/�/�/ �/�/����1?� X?j?|?�?�?�?�?�? �?�?OO0O�TOfO xO�O�O�O�O�O�O�O __,_>_�/?!?�_ E?�_�_�_�_�_oo (o:oLo^opo�oAO�o �o�o�o�o $6 HZl~�O_a_s_ ��_�� �2�D�V� h�z�������ԏ�o �
��.�@�R�d�v� ��������П⟡� �'��N�`�r����� ����̯ޯ���&� 8�I�\�n��������� ȿڿ����"�4�� U��y�;��ϲ����� ������0�B�T�f� xߊ�I����������� ��,�>�P�b�t�� Eϧ�i���Ϗ��� (�:�L�^�p������� �������� $6 HZl~���� ������/��V hz������ �
//./��R/d/v/ �/�/�/�/�/�/�/? ?*?�3W?�?C �?�?�?�?�?OO&O 8OJO\OnO�O?/�O�O �O�O�O�O_"_4_F_ X_j_|_;?�?_?�_�_ �?�_oo0oBoTofo xo�o�o�o�o�o�O�o ,>Pbt� �����_�_�_�_ %��_L�^�p������� ��ʏ܏� ��$��o H�Z�l�~�������Ɵ ؟���� �2��� �w�9�����¯ԯ� ��
��.�@�R�d�v� 5�������п���� �*�<�N�`�rτ�C� U�g��ϋ�����&� 8�J�\�n߀ߒߤ߶� �߇������"�4�F� X�j�|�������� ��������B�T�f� x��������������� ,=�Pbt� ������ (��I�m/��� ���� //$/6/ H/Z/l/~/=�/�/�/ �/�/�/? ?2?D?V? h?z?9�?]�?��? �?
OO.O@OROdOvO �O�O�O�O�O�/�O_ _*_<_N_`_r_�_�_ �_�_�_�?�_�?o#o �OJo\ono�o�o�o�o �o�o�o�o"�OF Xj|����� �����_'ooK� u�7o������ҏ��� ��,�>�P�b�t�3 ������Ο����� (�:�L�^�p�/�y�S� ��ǯ��� ��$�6� H�Z�l�~�������ƿ ������ �2�D�V� h�zόϞϰ��ρ��� �����ۯ@�R�d�v� �ߚ߬߾�������� �׿<�N�`�r��� �����������&� ����	�k�-ߒ����� ��������"4F Xj)����� ��0BTf x7�I�[����� //,/>/P/b/t/�/ �/�/�/{�/�/?? (?:?L?^?p?�?�?�? �?�?��?�O�6O HOZOlO~O�O�O�O�O �O�O�O_ _1OD_V_ h_z_�_�_�_�_�_�_ �_
oo�?=o�?ao#O �o�o�o�o�o�o�o *<N`r1_� �������&� 8�J�\�n�-o��Qo�� uow�����"�4�F� X�j�|�������ğ� �����0�B�T�f� x����������ᯣ� ��۟>�P�b�t��� ������ο���� ՟:�L�^�pςϔϦ� �������� ��ѯ� ��?�i�+��ߢߴ��� ������� �2�D�V� h�'ό��������� ��
��.�@�R�d�#� m�Gߑ���}����� *<N`r�� ��y���& 8J\n���� u�������/��4/F/ X/j/|/�/�/�/�/�/ �/�/?�0?B?T?f? x?�?�?�?�?�?�?�? OO���_O!/�O �O�O�O�O�O�O__ (_:_L_^_?�_�_�_ �_�_�_�_ oo$o6o HoZolo+O=OOO�osO �o�o�o 2DV hz���o_�� �
��.�@�R�d�v� ��������}oߏ�o� �o*�<�N�`�r����� ����̟ޟ���%� 8�J�\�n��������� ȯگ����Ϗ1�� U��|�������Ŀֿ �����0�B�T�f� %��ϜϮ��������� ��,�>�P�b�!��� E���i�k������� (�:�L�^�p���� ��w����� ��$�6� H�Z�l�~�������s� ��������2DV hz������ �
��.@Rdv �������/ ����3/]/�/�/ �/�/�/�/�/??&? 8?J?\?�?�?�?�? �?�?�?�?O"O4OFO XO/a/;/�O�Oq/�O �O�O__0_B_T_f_ x_�_�_�_m?�_�_�_ oo,o>oPoboto�o �o�oiO{O�O�O�O (:L^p��� ���� ��_$�6� H�Z�l�~�������Ə ؏�����o�o�oS� z�������ԟ� ��
��.�@�R��v� ��������Я���� �*�<�N�`��1�C� ��g�̿޿���&� 8�J�\�nπϒϤ�c� ���������"�4�F� X�j�|ߎߠ߲�q��� ���߹��0�B�T�f� x������������ ��,�>�P�b�t��� �������������� %��I�p��� ���� $6 HZ�~���� ���/ /2/D/V/ w/9�/]_/�/�/ �/
??.?@?R?d?v? �?�?�?k�?�?�?O O*O<ONO`OrO�O�O �Og/�O�/�O�O�?&_ 8_J_\_n_�_�_�_�_ �_�_�_�_�?"o4oFo Xojo|o�o�o�o�o�o �o�o�O_�O'Q_ x������� ��,�>�P�ot��� ������Ώ����� (�:�L�U/y��� eʟܟ� ��$�6� H�Z�l�~�����a�Ư د���� �2�D�V� h�z�����]�o����� �����.�@�R�d�v� �ϚϬϾ������ϳ� �*�<�N�`�r߄ߖ� �ߺ����������ӿ �G�	�n����� ���������"�4�F� �j�|����������� ����0BT� %�7�[����� ,>Pbt� �W�����// (/:/L/^/p/�/�/�/ e�/��/�?$?6? H?Z?l?~?�?�?�?�? �?�?�?? O2ODOVO hOzO�O�O�O�O�O�O �O�/_�/=_�/d_v_ �_�_�_�_�_�_�_o o*o<oNoOro�o�o �o�o�o�o�o& 8J	_k-_�Q_S �����"�4�F� X�j�|�����_oď֏ �����0�B�T�f� x�����[���� ���,�>�P�b�t��� ������ί�򯱏� (�:�L�^�p������� ��ʿܿ���џ� E��l�~ϐϢϴ��� ������� �2�D�� h�zߌߞ߰������� ��
��.�@���I�#� m��YϾ�������� �*�<�N�`�r����� Uߺ�������& 8J\n��Q�c� u�����"4F Xj|����� ���//0/B/T/f/ x/�/�/�/�/�/�/�/ ���;?�b?t?�? �?�?�?�?�?�?OO (O:O�^OpO�O�O�O �O�O�O�O __$_6_ H_??+?�_O?�_�_ �_�_�_o o2oDoVo hozo�oKO�o�o�o�o �o
.@Rdv ��Y_�}_��_� �*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n��������� ȟڟ쟫��1�� X�j�|�������į֯ �����0�B��f� x���������ҿ��� ��,�>���_�!��� E�Gϼ��������� (�:�L�^�p߂ߔ�S� �������� ��$�6� H�Z�l�~��Oϱ�s� ������ �2�D�V� h�z������������� ��
.@Rdv ���������� ��9��`r�� �����//&/ 8/��\/n/�/�/�/�/ �/�/�/�/?"?4?� =a?�?M�?�?�? �?�?OO0OBOTOfO xO�OI/�O�O�O�O�O __,_>_P_b_t_�_ E?W?i?{?�_�?oo (o:oLo^opo�o�o�o �o�o�o�O $6 HZl~���� ���_�_�_/��_V� h�z�������ԏ� ��
��.��oR�d�v� ��������П���� �*�<������C� ����̯ޯ���&� 8�J�\�n���?����� ȿڿ����"�4�F� X�j�|ώ�M���q��� ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������ %���L�^�p������� �������� $6 ��Zl~���� ��� 2��S �w9�;���� �
//./@/R/d/v/ �/G�/�/�/�/�/? ?*?<?N?`?r?�?C �?g�?�?�/OO&O 8OJO\OnO�O�O�O�O �O�O�/�O_"_4_F_ X_j_|_�_�_�_�_�_ �?�?�?o-o�?Tofo xo�o�o�o�o�o�o�o ,�OPbt� �������� (��_1ooU��Ao�� ��ʏ܏� ��$�6� H�Z�l�~�=����Ɵ ؟���� �2�D�V� h�z�9�K�]�o�ѯ�� ��
��.�@�R�d�v� ��������п����� �*�<�N�`�rτϖ� �Ϻ����ϝ�����#� �J�\�n߀ߒߤ߶� ���������"��F� X�j�|�������� ������0����� u�7ߜ����������� ,>Pbt3� ������ (:L^p�A�� e����� //$/6/ H/Z/l/~/�/�/�/�/ �/��/? ?2?D?V? h?z?�?�?�?�?�?� �?�O�@OROdOvO �O�O�O�O�O�O�O_ _*_�/N_`_r_�_�_ �_�_�_�_�_oo&o �?Go	Oko-O/o�o�o �o�o�o�o"4F Xj|;_���� ����0�B�T�f� x�7o��[o��Ϗ��� ��,�>�P�b�t��� ������Ο���� (�:�L�^�p������� ��ʯ��ӏ����!�� H�Z�l�~�������ƿ ؿ���� �ߟD�V� h�zόϞϰ������� ��
��ۯ%���I�s� 5��߬߾�������� �*�<�N�`�r�1ϖ� �����������&� 8�J�\�n�-�?�Q�c� ��������"4F Xj|������ ��0BTf x��������� ��/��>/P/b/t/�/ �/�/�/�/�/�/?? �:?L?^?p?�?�?�? �?�?�?�? OO$O� �/iO+/�O�O�O�O �O�O�O_ _2_D_V_ h_'?y_�_�_�_�_�_ �_
oo.o@oRodovo 5O�oYO�o}O�o�o *<N`r�� ����o���&� 8�J�\�n��������� ȏ�o鏫o��o4�F� X�j�|�������ğ֟ ������B�T�f� x���������ү��� ��ُ;���_�!�#� ������ο���� (�:�L�^�p�/��Ϧ� �������� ��$�6� H�Z�l�+���O����� ������� �2�D�V� h�z��������� ��
��.�@�R�d�v� ��������}��ߡ��� ��<N`r�� ������� 8J\n���� ����/���� =/g/)�/�/�/�/�/ �/�/??0?B?T?f? %�?�?�?�?�?�?�? OO,O>OPObO!/3/ E/W/�O{/�O�O__ (_:_L_^_p_�_�_�_ �_w?�_�_ oo$o6o HoZolo~o�o�o�o�o �O�O�O�O2DV hz������ �
��_.�@�R�d�v� ��������Џ��� ��o�o�o]����� ����̟ޟ���&� 8�J�\��m������� ȯگ����"�4�F� X�j�)���M���q�ֿ �����0�B�T�f� xϊϜϮ���ѿ���� ��,�>�P�b�t߆� �ߪ߼�{��ߟ��ÿ (�:�L�^�p���� �������� ����6� H�Z�l�~��������� ��������/��S ������� �
.@Rd#� �������/ /*/</N/`/�/C �/�/{�/�/??&? 8?J?\?n?�?�?�?�? u�?�?�?O"O4OFO XOjO|O�O�O�Oq/�/ �/�O	_�/0_B_T_f_ x_�_�_�_�_�_�_�_ o�?,o>oPoboto�o �o�o�o�o�o�o�O _�O1[_��� ���� ��$�6� H�Z�o~�������Ə ؏���� �2�D�V� '9K��oԟ� ��
��.�@�R�d�v� ������k�Я���� �*�<�N�`�r����� ����y���������&� 8�J�\�nπϒϤ϶� �������Ͻ�"�4�F� X�j�|ߎߠ߲����� �����˿ݿ�Q�� x������������ ��,�>�P��a��� ������������ (:L^�A� e���� $6 HZl~���� ���/ /2/D/V/ h/z/�/�/�/o�/� �/�?.?@?R?d?v? �?�?�?�?�?�?�?O �*O<ONO`OrO�O�O �O�O�O�O�O_�/#_ �/G_	?_�_�_�_�_ �_�_�_�_o"o4oFo XoO|o�o�o�o�o�o �o�o0BT_ u7_��oo��� ��,�>�P�b�t��� ����ioΏ����� (�:�L�^�p������� e��ӟ���$�6� H�Z�l�~�������Ư د����� �2�D�V� h�z�������¿Կ� �����۟%�O��v� �ϚϬϾ�������� �*�<�N��r߄ߖ� �ߺ���������&� 8�J�	��-�?ϡ�c� ���������"�4�F� X�j�|�����_����� ����0BTf x���m�������$FMR2_�GRP 1Z��� ��C4  B��	� ��;M8E�� F@ cǂ5Wo�
8J���NJk�I'�PKHu��IP��sF!��{?ǀ  ��89��<9�8�96C'6<�,5��{Ag�  /+BH5�B�10 !@�3]3;"�33�7x]/n-8@UUT�*�@9 � {��>u.��>*��<����{>���>���l=<��=��U�=�v!>1�
{:�ܜ:�2B8'Ŭ9�IR7���9f�͛/$?o/!?Z?�E?~?i?�?��_C�FG [T ��?�? OO�;N�O 
F�0HA M@�<RM_�CHKTYP  ���&(� R{OMc@_MINi@������@�T X�SSB�3\�? 9�O���C�O�O�5TP__DEF_Oz���&	WIRCOM�h@_�$GENO�VRD_DO�F���G]THR�F dzdUdMT_ENB9_{ MPRAVCu]�G�@ �[�F@ G��@�GAw\H͊#Iv0�Iά �?�Oo�o(oK*� �QOUc�PAKRK<�@��oIo�o�o��o��C�  D��o�h1A|A$ B��L.rN�i�O�PSMTd�Y*�@t�$HOSTC�2s1e�@����7 MC��T{����  27�.02�1�  e�_�q�������M��Ə؏��������	�anonymous#�Q�c�u��������6������� F�'�9�K�]�o����� ����ɯ쟆�0��#� 5�G�Y�k�����ҟ�� �׿�����1��� �g�yϋϝ������ ����	��-�p��ϔ� ���ߺ�ܿ�������� �H�)�;�M�_�q�� ���Ϲ��������D� V�h�z�|�R��ߑ��� ���������!3 Eh������� ��*�<�N�PA�� ew������� �//<n3/a/s/ �/�/�/���/$/ ?X9?K?]?o?�?� �?�?�?�?�/�?B/#O 5OGOYOkO}O�/�/�/ �O�?�O,?__1_C_ �?g_y_�_�_�_�OT_ O�_	oo-o?o�~�q�ENT 1f�y��  P!�_�o  �p~o�o�o�o �o�o'�o3\ �D�h���� ���G�
�k�.��� R���v���鏬��Џ 1��U��N���z��� r�ӟ�������ޟ,� Q��u�8���\����� ᯤ����گ;���_��"�QUICC0 l�H�Z���~�1�������~�2����[��!ROUTER�\�8�Jϫ�!PC�JOG�χ�!�192.168.�0.10��z�CA�MPRT����!b��1��#�
�RTu��'�9ߚ� !So�ftware O�perator Panelw������`dNAME !~mj!ROBO����S_CFG 1�emi ��Auto-st�arted�DFTP�O���O�_�� �O��������c_>� P�b�t����+����� �����@\�n�� a����x���� ��'9Kn� �������O�O �O�OV,/�k/}/�/ �/�/v�/�/�/?? B/�/U?g?y?�?�?�? �//(/*?O^/?O QOcOuO�OJ?�O�O�O �O�OO�O)_;_M___ q_�_�?�?�?�_�O�_ 2Oo%o7oIo[o_o �o�o�o�_�olo�o !3EW�_�_�_� �o�o�����o A�S�e�w����.��� я�����\n� �s��������͟ߟ 񟴏�'�9�K�]��� �������ɯۯ�0� B�T�f�h�Y���}��� ����ſ������� 1�T�ֿg�yϋϝϯ������_ERR �g�����PDUS_IZ  V�^t�����>	�WRD� ?J�7�� � guestV�I�[�m�ߑߣ����SCDMNGR�P 2hJ����7�V�8V��K�� 	P01�.03 8� �  e�?���  ;  ��  � ��������@��-�������x����0���y� d����,�>�P������  	D��d����������_GROU��i*������	���]5{�QUP�3��������TYC �����TTP_A�UTH 1j��� <!iPen'dan��%`Ϗ��!KAREL�:*%.@KC�UewM VISION SET����V�K�� J(@:�^p�����CTRL� k����%V�
�4�FFF9�E3�5�FRS�:DEFAULT�3,FANUC� Web Server3*! 5���1� C���/�/�/�/�/?���WR_CONF�IG l�� �3/��IDL_C_PU_PCR V�sB�8�u0 BH[5�MINf<!�y5GNR_IO���V����]0NPT_SIM�_DO�6�;STAL_SCRN�6� ���INTPM?ODNTOL�7�;�!RTY�8u1�6� N��ENB�7��Y4OLNK 1m��E�}O�O�O�O�O�O|�OaBMASTE�0���aBSLAVE �n��URAMCOACHE_�2O��O_CFGI_`CaS�UO��l_]RCMT�_OPR �2�ʟSY�CLH_{UL _AS�G 1o��#�
 �Oo o2oDoVoho zo�o�o�o�o�o�o�o\�K�RNUM����
]RIPF_XWRTRY_CN�_{U�1(���|A��� ]R�PfRp'^=з=�]0�P_MEMBER�S 2q��� $�%�r����w���]0RCA_AC�C 2r��  �V�

 O��V�6IP_��s"S�d�^�h�Z���28��BUF001 2�s��= 	�u0  u0	�քU�ք�ք�ք�ք��փ

�7��  7��փ����փ.��.�#.�2.�D.�S�.�d.�t.��.���.��.��.��.��j.��.��փ��U��(��8��I���X��j��yփ �"��"�� ��0�A�P�b��q���������քքք&�ք5քFքVքgJքvք�փ��2�� ҃ց܁����� �������ց�� ���ց$�)�-�ց 4�9�=�9�E�9�M�9� U�9�]�9�e�9�m�9� u�9�}�9���9���9� ��9���9���9���ց ��������Ő��͐�� Ր��ݐ��吹��ց �������������� ������%���-��� 5���=���E���M��� U���]���e���m�� u��}�ᢅ�ᢍ�� ��ᢝ�ᢥ�᢭����ց��3ɯ҅�� ��������� "�#�*�%�3�&�4� C�B�E�S�B�U�c�B� e�s�B�u���B҅��� Bҕ���Bҥ���&� ó��Œӳ��Ւ��� ��&������� ��#��%�3��5� C��E�S��U�c�� e�s�U�u���U򅢓� U򕢣�U򥢳�U�,��gQ2t��4,%��&�<&�K���2�5�HIS��v��� �S� 2023-07-19Y& |B;�_�l� ~���������������^V�sE�8Q� J\n���W'��Y!׀������s!�^��s  77��q5" 4FXj|��� ���//0/B/ T/f/x/�/�/���/ �/�/??,?>?P?b? t?�/�/�?�?�?�?�? OO(O:OLO�?�?�? �O�O�O�O�O�O __ $_~#�Ƞ/�A�S�j�dU��R3_�_�_�_�_ �_�_o!o!3io�{o�o�o�o�o�� �c� �^� �b� -�  L� 8  ^iO{OASew ������eO, �+�=�O�a�s����� ������ȏ��'� 9�K�]�o�����ʏ܏ �۟����#�5�G� Y�k�}���Ɵ��ůׯ �����1�C�U����T_f_S�ө��� ȿڿ����"�4�F� 4oFoXo�Ϡϲ����� ���oQ����Q�� Q�� ������j�|ߎ� �߲����������C� U�B�T�f�x���� �������-��,�>� P�b�t����������� ���(:L^ p����������  $6HZlZ��l�I_CFG 2�wz� H
C�ycle Tim}e�Busy��Idl��m�in}�U�p��Read>�Dow��� ��Cou�nt�	Num D����`,w�7!�EQPROG�xz����p/�/�/��/�/�/?�@USD�T_ISOLC � z��pJ�23_DSP_ENB  B;�c0?INC ys=w��P0A   ?� � =���<#��
O1�9:�o ��1�?�?���?	O]6OB� Cl3��6"A�G_GROUP �1zB;�b<A� �3�	nOO?��/�Ow�Q�O�O�O�_�O0_B_T_f_���?IG_IN_A�UTO/D�:c0PO�SRE*O<FKANJI_MASK�V��ZKARELMO�N {z�h/w�y +_DoVohozo�o�bJ�#|�'~3w��e|�_4KCL_L�P�NUMp0�o$KE�YLOGGING��`��bA{5� LA�NGUAGE �z�Jp�DEFAULT Xq6h�LG�}�*���w�x�0�  }v�H  �w��'0��w��w��?)7;��
�q(?UT1:\�o� ����0�=�@O�a�x�������(3o��c�LN_DISP ~�?��O�O>��OCTOL9�w��Dz� K1�1O�GB'OOKq0i}d���������X�|���� ϟ����us�'��	m��yjA%;o��?�1k�_BUFFw 2�B; �w�2�����*2ү� � �-�$�6�c�Z�l� ������Ͽƿؿ����)� �2�_π3��DCS ��)�2�1$� c�����������v��IO 2��� 1�3�jA�6�F� X�j�~ߎߠ߲����� ������0�B�V�f� x����������տER_ITM?>d �_?�Q�c�u������� ��������); M_q���I��SEV�`s=�TYP?>.�!3���QRSTt�S�CRN_FL 2��� ��ϧ�����//DTP�p??�C�NGN�AMl4��Jrr�UPMS�GI\�U{5}�!_LOAD'@�G %@*%D�MAYɥ�/G�MA?XUALRM�b�Q�C��{5
�"�!_PR�$�P a�%�� C��i�ٯè�)3H@P 2�w�k �Ʀ	O!t�0��0�P?���2�?�? �?�?���?+OOOO2O DO�OpO�O�O�O�O�O _�O'_
__]_H_�_ l_�_�_�_�_�_�_�_ �_5o oYoDo}o�oro �o�o�o�o�o�o1 UgJ�v�� ���	��-�?�"� c�N���j�|������ ̏����;�&�_�B� T���������ݟ�ҟ����7��'DBGDEF �25?1>1�@�R�_LDXDI�SAm ?+�MEM�O_APg E ?=@+
 d�� ��ү�����,�>��� FRQ_CFG� �27h�A ��@���!�<?4dA%A���R�d�z2�2;��4*z��/�� **:� !���ȟ�!�,�>�k� b�tϡϘϪ���#�25� �����'�� �6�,(��~���lߩߐ��� �������'��K�]� D��h�������*?ISC 1�@)� �)�#��4i�9�$��r�]�������_MS�TR ����S_CD 1������ ��,P;t_ q������ &L7p[� �����/�6/ !/Z/E/~/i/�/�/�/ �/�/�/�/ ??D?/? A?z?e?�?�?�?�?�? �?�?OO@O+OdOOO �OsO�O�O�O�O�O_ �O*__N_9_^_�_o_ �_�_�_�_�_�_o��MKg������&o$MLTARMf���۷Qb ��b��o�dQ�METsPU��b�����NDSP_ADC�OL�ef��nCMNmT�o �eFN�`|�o�gFSTLIw�� ���g~�c��t�ePOSC�F5w�nPRPMl�o�yST�`1���w 4��#�
� ���!��!�#�5� w�Y�k��������ŏ ׏����O�1�C����o��aSING_C�HK  $M7ODAe���Ok�Qn��DEV 	���	MC:�HOSIZE��`ȿ�TASK %���%$123456�789 `�r���T�RIG 1��� lQ�����Lٮ�﯌L�B�YP-�L�Ք���EM_INF �1�ۻ`)�AT&FV0E0���k�)S�E0V�1&A3&B1&�D2&S0&C1�S0=Z�)ATZk�����Hÿ�z�߯Ϣ�A�C���g�Nϋϝ� Q���u��� �����Ͽ@�w�d�v� )Ϛ�U߾��߷��ߧ� ��*������r�}�7� �����������&� �J�\���3�E�W� i�������5�4�� X|�u�e�w� �������0B��f ��EO�{�� //�>/�' �/K�/�//�/�?��/'?L?3?p?�NIwTORPpG ?��   	EX�EC1c�22�83��84�85�8���67*�88�89c�2:" D�2D�2D�2D�2 D�2D�2D BDB�DBC2%H21H2�=H2IH2UH2aH2�mH2yH2�H2�H3�%H31H3�2��R_�GRP_SV 1ݔ@� (w����<� ��>%���6���?�u=���J��_D20�ySION�_DBɐ�͝a�  �p�p�放U��p��W��  
v�f0N �  E��P��[��`�P�-ud�1�/oAoSo�aPL�_NAME !�Q�|`�!De�fault Pe�rsonalit�y (from �FD)�P�bRR2�7Q 1�L�X�L�x|a�P dzr�o�o�o�o #5GYk}�� �������1�C���2�on����������ȏڏ������< ]�:�L�^�p����������ʟܟ� �[i*�D)�:�
)�^�]dPM� ��������ү���� �,�>�P�b�t����� g�y�ο����(� :�L�^�pςϔϦϸ� ���ϫ����$�6�H� Z�l�~ߐߢߴ����������� �2� �F@ G&h �G��]gSP  �_�q�]bd[�C��� �������D�7�Zj���	���=�@�  -�X�N�`�r�������@��SP�0��	]b-��	`B�<N`:�oA�b���~� A�  �	�W�V]`�S �]`��PCT��s�  h��)�  �  u$ �T&"�C�gydН��\kR6R 1�ti�P*0 �� f2|`  �@D�  !?�>#X,?]`!]aA/��%�XJ.�;�	l,"	 ���pJ�n �NP`e  Կ � � �� �� ��"SPK��K ��K=*��J���J���J9٧�U�p��/SP@_f��"j?�@�(E14!��/�#�N�����;f,1�� �a_������-�@o¾  T1�HZ0�Z0� �/  >c��=��>�]a������l? �?�2-!�3�&�. p�Pm P�� ��P�  ���P�F�*O�%	'�� � HBI�� �  ����&:�ÈlOß�=��̈́E�"@�O�@�>!�O/K"��&&�&�Q_�  '.T�!-0@2��@����"Z=0@A?C� C�P_C�� Ca0Ce0uCi=%��A�%� 0 �P�l�-hhX�'B�P�Q���A�U]aDz�on?3oo Coio�O�dIA�R�TZ�v�A���  �4@?�ff���o�o�no  #{�!8�@9Gz>L�@�0(!�*(�@uu�0�v�i{!Ht#t$�C?]t�@,���<
6b<߈�;܍�<�ê�<���<�^�Ȭ/�C�A�K"��#,"� ?fff?�@?&&���@�.�8��J<?�\�D�N\��I�R!� -$�)%|�'��
�`$ �oЏ���ߏ��<��'�`�r�]����He�FiP��ҟ����m����J��F�  �F���BG�d GC�qV���R���ů ���ԯ���1��U� @��O���F�IG/�ӿ 1���m��0�B�T�:�9��o�{�33ϩπ��ϸ������{An� ��_�EC��U���<��d�?�؃ߊ�h�߮��I�i4����C CfPa0�¸�Ԑ0؜�@�@I����B>�)A��C�AIA���@�?�\������@ �������=q�A��Ay�I�33@0��@���C�1�������(��Cb��=q��Ů�����H�� G��� G�B�I��(E�� C�e��� I"L�J��HV@G5� E�x C���I3�J0��G���I�� 0 C='�߀�k��� ������������" F1jUg��� ����0B- fQ�u���� �/�,//P/;/t/ _/�/�/�/�/�/�/�/ ??:?%?7?p?[?�? ?�?�?�?�? OO�? 6O!OZOEO~OiO�O�O �O�O�O�O�O __D_ /_h_z_e_�_�_�_�_t�_y�(������r��$e�U���o&o9�3�8�x@oRo9�4Mgulo<~o9ѴVwQ�o�o�4p�+4�] �m�i�o(L:|Ju�P�rP~~�������_�����{R��G�2�W�}�h�  �`��ˏ�� �ڏ����F�4�j�X�p�z��������ԟz����4�"��X�F�|���  2 �F@9�G&h6����9�B�&��L)��C�&�9�@-� �9�o�+�=�O���� ���Ħ�GA�w\]�����ɿ7�?Q��|p9�t�9��9���{�
 ֿ9�K�]�oρϓ� �Ϸ����������#��z����hk�y���$MR_CA�BLE 2�hxO �ћqT�p@����?>𦡆і����кƠ��C���ޱO8�tB�=�;�m�or�ް�F
޶�ߕ���>��š��C�N��|�����a^��vްޱE�Cx�e����L  ����C֠:���:���▋(ްO�N����"�4��ՠ��y�By�ԡ��HE鈢�lt�޵;5�~v�/ߘ���k���� ��C��L�>�8�f�\� n�������������?(��H�� oq<� ��ܸ���ܸw*,** \��OM �i�������Ӫ�%%� 2345678'901i{ f�D�ް�ް�!�ޱ�
�not? sent 5��WpuTES�TFECSALG&#�egۺ�d.$�0����ы��p���޷Y/k/}/�/ 9�UD1:\ma�intenanc?es.xml�/�/�  ��D?EFAULTa�\ҿGRP 2�M � pė�޵  ��%1st m�echanical check�ޱ�z3鰄1�?��[ph��?�?�?�?��?޲R3controllerb4,O{?PO���?|O�O�O�O��OAMY=�O޲"�8SްQ_���kG8_J_\_n_�_�JC O�__�_�6/_o�o(o:oLoBC[0g�eW2. batt�eryPo�_�o��	 �_�o�o�o�o_i@�dui@able  D50Pq����`���o������AddgreaYs;޷f��-ް�#���{P�b�t�h����A
ddoi�/��+�?��&�8�J�\�Adj7޶����<ް������
�؟���� �#|!too�����>ǟ��ய��ү�AOv�erhau�Ow��"� xް,�3�:5��`�r�������ްA$Q�пSV�� O� $�6�H�Z�lϻ���߿ �Ϲ������ �2� ��VߥϷ��Ϟ߰��� ����5ߝ��k��� d�v���������� 1��U�*�<�N�`�r� ������������ &8��\����� �������M" q�X�|��� ��7I/mB/ T/f/x/�/��/�/ �/3/??,?>?P?�/ t?�/�/�/�?�?�?�? OOe?:O�?�?�?�O �O�O�O�OO�O _OO �OsOH_Z_l_~_�_�O �_�__�_9_o o2o DoVo�_zo�_�_�o�_ �o�o�o
ko@�o �ov�o����� 1�Ug<��`�r� �������̏�-�� Q�&�8�J�\�n����� ��ȟ�����"� 4���X�����˟���� į֯���I��m�� ��f�x���������5��	 T¿��� *�4�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ߮��� ��������,�>�P��b�t����� � �b�?�  @�  ���	������H�Z�l��*��** @�>�7� ����������,>��e�^���A ���u���E Wi�Ugy�� ���/�/-/ ?/�/u/�/�/�� /�/�/??�/;?M?�_?�/�/���$�MR_HIST �2�>��0� 
� \
�$ 2345678901�?(�4�?���?9�)O ;O�?$O��O�O�O^O pO�O�O_�O�O_I_ [___6_�_�_l_�_ �_�_o�_3o�_Woio  o�oDo�o�ozo�o�o��oA�d�0SK�CFMAP  .>��08�1��`IYuONR�EL  �5�rq�0[rEXCFE�NB�w
psXu�qF�NC��tJOGO/VLIM�wd�3��[rKEY�w��_PAN�x+�'��[rRUN �,�SFSPDTYP�x<�uZsSIGN��t�T1MOT��q�[r_CE_GRP7 1�>�rs�2 ڰ9���c��8��8&� g����B�����x�� ��ڟ�ҟ?�Q��u� ,�����b�ϯ��ȯ� ��)�;�"�_�������|����7[qQZ_E�DIT��lw��TC�OM_CFG 1��h}�u�&�8� }
��_ARC_�r��5�yT_MN_oMODE����yUAP_CPL]���tNOCHECK� ?h{ @ ��������,� >�P�b�t߆ߘߪ߼�����ߍ{NO_WA�IT_L���ՀN�T���h{w��c�2�_ERR߁2�hy�1�6�����*���q�����w�O`�>g�| O����0�r�a<O�00 ?�5��O�5��p"�Y�PAR�AMa�h{���� ������1�� = O08Z lHx���������.��R~��ODRDSP\�����xOFFSET�_CAR�bψDsIS��S_Aw��ARK���OPE?N_FILE����;��S�OPTIO�N_IO!�3� M_PRG %hz�%$*E/W.�WO������p00�%�d.2  p��v� C�!	 ч�h�!�f����hRG_DSBL'  �7rqK�?�eRIENTTO��p�aC��pqqA� fUT_SIM�_D'or��hV~lLCT �<�粛$;��9�ed`7_�PEX���4RA-T� d�u�4��UP �q>��{ �OOOBOPI��$��2ރ�L��XL�x[3�0C�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o�g2�O/oAoSoeowo �o�o�o�o�oB�o�o 1CUgy� ������f�o�~9@�!�N�P�K�]� o���������ɏۏ� ���#�5�G�Y�(�:� ������şן���� �1�C�U�g�y����� l�~�ӯ���	��-� ?�Q�c�u���������`Ͽ�s�¯��� � 2͠4A�!S�e�Gυ� ����A�����ϭ�������!�3�Q� W�uߗ���{ ��������	`����!�x�:�o@1?�Q�c�|u�A�  ��
V+��!+�21� �9���s  �h�p )  ?�  u$�� ���)��&�_�J����^fBl@O�01� �� � {D}��0 ��$�  �� @D�  ���?���X,q?+���+�D��������  ;�	�l��	 �߀pJ3 ������*  � � w� �I � �O�u�H(��H3k�7HSM5G�2�2G���GNɁ3h��(ϙ�u�C)H50�R50������r�û�¾  ��� �� �)���m�AK�µ�+�²���801 io���u����� p m�3�P00� �  � ��u��q�	'� � "�I� �  ����o�=���81/C+�@Y/_  Z�!�/��"������q�NA0�/  '�R0�$���CA0C�	��*C. ??�q��p�Az
b0�lwhhXn�B� �1��~�p!�5��zn��?3�?�?O .OU/GD!N2K4a+�Ӻ���@?��ff�ϏO�O3O !���O�KA8+��O�Z>LS ���J( +�:U�EV^I@99ң#?"T� ,A<
�6b<߈;����<�ê<�?��<�^�q�_2�AAp+���#���?fff?p ?y&�PD@�.�R�J<?�\�	bN\��U2�Q�@ ��Ao��`o�W%�O�o �o�o�o�o�o�o% 7"[mD�|��,oNoPo���xF��  F��+�G�d GCFQ�T�� d���u�����ҏ���� ����/M��&
 ������2�����d��J��O�[�3p ޟw�b�������
<�!A3�墚?+�C���x��w�)�?��H��O���s�
�4����C��C�࿇��b��b�a��@I��	B>�)A��C�AIA���@�?�\��������@ �������=q+�R!>�I�33@0��@���C�1����[�����C'��=q��Ů���	H�� G��� G�B�I��(E�� C�^l���I"L�J��HV@G5� E�x C����I3�J0��G���I�� E@� C��E� 0�i�Tߍߟߊ��߮� �������/��,�e� P��t�������� ���+��O�:�s�^� ��������������  9$]oZ�~ �������5  YD}h��� ����/
/C/./ g/R/d/�/�/�/�/�/ �/	?�/-???*?c?N?Ї?r?�?>�(I��ٙ^opR���5�5����?�?@�3��8�OO@�4Mg�u1OCO@��VwQ�]OoO4p�+4�]�M�I�O�O�O�O(_�L:�P�RPC^>�_�l_�?x_�_�_�_�[R�_�_o�_o,Bo-o  �@�EoWo �o{o�o�o�o_Q��o/{5?u c���?��������A�O�  �2 F@@�G�&hl���@�B�0���ձC��@�@򯷏ɏۏ����"�@��oL�^�p������@�?���AP@�J�d@�@�<���@�
 �����"� 4�F�X�j�|�������`į֯�?ʶ���-K��y��$PA�RAM_MENU� ?�E��  DEFPULSE���	WAITTM�OUTL�RCV�_� SHEL�L_WRK.$CUR_STYLJ�;��OPT�����PTB����C��R?_DECSNW�4U ���%�N�I�[�m� �ϑϣϵ����������&�!�SSREL_�ID  �E]Q��5�USE_PRO/G %0�%"߇�6�CCRc�G�]Q8����_HOST �!0�!���ߔ�T TP���ӿ�����4�>��_TIMEa�G����!�GDEBU�GE�0�6�GINP?_FLMSK]��qT�P���PGA��e |�;���CH��^��TYPE-�9�!��Q�z�u����� ��������
) RM_q���� ���*%7I rm������/��WORD ?�	0�
 	PyRy��SMAI����RSUͱ=#TE���S�	��J"CCOL�Uf)�/��LcЫ �@��`ȯ�d�q�TRACECToL 1��E:�� AP� ��'AP;P�.�&DT� Q��E0� �D � � ���[Q12�� 12Ԑ12��12̐12Ȑ�10� _4_4�_4G�10� 4�444���2_463�=4�E4�!`3�V3�54�=4�E4��M4��6^5^5_4*_4	_4
_4_4.?@@?R?d?v?�?�9�DT�A@�ED�MD�UDU�]D�eD�ED�MD��UD�]D��FnC�TVC�D�%D�-DU�5D�=D�ED�MDU�UD�]D�eD�V�vC�}D��D��D�K �D�D�E�O �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�o �o�o1CUg y�������dU�d�d �d!�d�"�d#�d$waN� ke'1[�o����� ����ɟ۟����#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� �ߧ߹��������� %�7�I�[�m���� �����������!�3� E�W�i�{�����k��� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�/ �/�/�/�/�/�/?? +?=?O?a?s?�?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O_#_5_G_Y_ k_}_�_�_�_�_�_�� �_oo1oCoUogoyo �o�o�o�o�o�o�o	 -?Qcu�� �������)� ;�M�_�q��������� ˏݏ���%�7�I� [�m��������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�e�w��� ������ѿ������#��$PGTRA�CELEN  �"�  ���!��7�_UP ����f��n�R�g�7�_�CFG �f��P�!�g�����ĭϸ�I���  ����{�DEFS_PD ��� ��I��7�H_CONFIG �fŮN� !�!�d�-��F�  �0�P�����L�!��7�I�N~�TRL �d�ͦ�8��a�PE�;���f��ĸ,Ѹ�7�LIDù���	��LLB 1}�� �M��B<�B4�� �M�%��Pպ� �<< �?� O�n�O�f����� �����"���<�j�P�r�����8����� ��
Q�@3Ev~��GRP 1�����"�@��
����!�AM��D�@ D�@ kCf� @ �1�`���	�	,�,����0uG���´F(BIpP:L��p�!�>�l7>�����/.� �=�-=%�T /Q//N/�/r/�/�/�0/�/�/�/?)?? G DzN3W?!�
>? ?.?�?�?�?�?�?�? �?!OOEO0OBO{OfOПO�O�O�J)�A
�V7.10bet�a1�� A�{�� R�!�A!���@?!G�Q=y��#�B���$Q@w����B�l�4Q@�A���QT �Oi_{_�_�_FTp���<��_�_�_ �_.� ��O��O�0o�Bo,ofoPo�o�A-�p��u0�mf��o� �o���@�AWP�R6�c B��B�>0uSBHfs�d!�!��PuM���d����r�cx�tx�����$|��� �0��<�-�@�F�0�A�33`��������KNOW_M  �"�����SV ��C�]�m? � �$��oH�3�E�~�!�����M��� ՔR	��ѐl�b��^���hhXd��1q� (�`0u8�4�����MR�³��&�oj3�������OADBANF�WD����ST�1� 1�f��4 �խY�!

��.�_� R�d�v��������п �'���]�<�Nϓπrτ��ϨϺ����2p����	�ݠ�<3���3�/�A�S��A4p߂ߔߦ��5���������6�(�:�L��7i�{�����8���������MA�֠��b�OV_LD  ���~�PARNUM�  �������S[CHa� o�
��p��	�UPD����#bb�_CMPa_��d����'�~zER_CHK����˒����RSu�ٯ��_MO�֯�_�a�_REWS_G����
V_ ��ch����� ��/
/;/./_/R/d/7�DT�/9 oУ/�/�/;���/? ?;�!?@?E?;h� `??�?;���?�?�?�;��?�?O;V �1��vߠ��@`�}\�THR_ICNRu�f��dqFoMASS~O Z�G�MN}O�CMON_�QUEUE �P���
�Qa�N �U�N�F�H SENqDQ#YEXE._�UD BE-P_ SO�PTIOW,PP�ROGRAM %�J%P<O��R?TASK_Ic�u^OCFG ��Ox���_
`DATA��M�kP�
2ʕ yo�o�o�o�olo�o�o 	-�oQcu�^:oINFO���Wm��DC����(� :�L�^�p��������� ʏ܏� ��$�6�H�4�w�t�Wl r)	a6��K_a�i�~��ENBd�ѹ�i2ԘGa2̙� X,		��=��� ���@	�N�9�$��8�8��`D��_EDIT ��o����dWE�RFLOXdC�RG�ADJ �}�A	����?
���AϦ�Q������?�  Bz��"ga<8�
�v%$�\�0èr-�g�2���rk	H�@locB{BP���q@'��ǽ*۰/ݲ **:�ֿ��qy��.@A��ſ��K�@�c���\I)#Ⱥ��1�[ϩ�g�������w�A.@u��� ����O���K�5�/�A� ��e߷ߡߛ߭�'��� #�����=��y� s������������� k��g�Q�K�]����� ��������C��?) #5�Y���� ���1 �mgy���� ��_/	/[/E/?/Q/ �/u/�/�/�/�/7?�/ 3???)?�?M?�?�?�?�?{�	&o0OŠO<WOBD�t$ qO�K�EO�OAO�O�O	�PR�EF ��Š�Š
ϥIORIT�Y�W���ӡMPD�SP�Q��A�7WUT��V��ΦODUCT��Q}��O��OGg�_TG���R���vRHIBIT_D�O���[TOENT� 1�}� (!AF_INEaP�og!tcp|oGm!ud6o~on!icm^o��vRXY��}��š)� ��o�oŠ��o�e�o: !^EW�{��������6�H�*uS���A�J�����^£>Ԥ�Ѷ�!/��z��¤�r�}��A;�,  � P}�8�J�\�n�ť�߆Zߏ����ҟ��£]�ENHAN�CE �i�}�A��dޏD�+�rV�D�� _SɡӡPOR_T_NUMbSŠ�.Uӡ_CAR�TRE���l	�S�KSTAaW�[SL�GS`ٸk��;�HPUnothingL�)�;�M�]����������_�TEMP څY���5�q�_a_seiban�OϯO(�N� 9�r�]ϖρϺϥ��� �������8�#�\�G� ��kߐ߶ߡ������� ��"��F�1�C�|�g� ������������� 	�B�-�f�Q���u��� ����������, P;`�q����������VE�RSI@P�WQ �disabl�e^���SAVE �ۅZ	267_0H769'��!4���po� !		(kR�?;+2/ES�eO/x/�/�/�/�*�g,��/z�n_�P +1ܸk�20
B�5<?N?�7�@URG�E�B�P�^�aWF z0�QdT�pVW`�4�LQ��WRUP_DELAY ݼ���5R_HOT �%FnQ3�O�5R_?NORMAL�8�Rx
O_O.GSEMI>O�dO�O�AQSKIP3�p�+3x�O __0_�M�5W_eWO_ �_�_�_o_�_�_�_o o'o�_Ko9ooo�o�o Yo�o�o�o�o�o�o 5#Ek}�U� ������1���U�g�y��5�$RB�TIF�4��RCV�TMOUէå]���DCR3��I� ��AC��}�C�&�C����?���>��9�<?��M���`�B	1��$,���"��@�N�OC�?_ �<
6b<���;܍�>u.��>*��<����U���?����� ��ߟ���'�9��K�]�o��������ER�DIO_TYPE�  !=����ED�PROT_CFG� ��G�4B�H3E���A2�n� ���B� � T�b�����:�����п ��c�ϐO(�G_I�;� Y�[�mϣϑ��ϵ��� ���ߡ���E�3�i� Wߍ�{ߝߟ߱���	� �-�/���?�e�S�� w������������ +���O�=�s�a����� ������������� K9o]����� ����5#E GY�}���� �/�1//U/C/y/�g/�/���/����I�NT 2��9J��ǱG;� ?&;s�x��N?�f�0 l? ~;�/�?�/�?�?�?�? �?OO,ORO@OvOdO �O�O�O�O�O�O�O_ *__N_<_r_`_�_�_ �_�_�_�_�_o&oo Jo8ono\o~o�o�o�o��o�o��EFPOS�1 1�̩  x�/:y�A?c N��x-?y�� ��"��F��C�|� ���;�ď_������ ���B�-�f����%� ��I��������,� ǟP�b����I����� ίi�򯍯����L� �p����/���ʿe� w������6�ѿZ��� ~��{ϴ�O���s��� �� �2������z�e� ��9���]��߁���� ��@���d��߈��5� G���������*��� N���K������C��� g���������J5 n	�-�Q�� ��4�Xj Q���q�� /�/T/�x//�/ 7/�/�/m//�/?? >?�/b?�/�?!?�?�? W?�?{?O�?(O:O�? �?!O�OmO�OAO�OeO��O�O�O$_�Cu2 1��O�O_�_{_ �_�O�_s_�_�_�_2o �_Vo�_zoo�o9oKo ]o�o�o�o�o@�o d�oa�5�Y� }�����`�K� �����C�̏g�ɏ� ��&���J��n�	�� -�g�ȟ��쟇���� 4�ϟ1�j����)��� M�֯q�����ϯ0�� T��x����7���ҿ m�����ϵ�>�ٿ� ��7Ϙσϼ�W���{� ߟ��:���^��ς� ߦ�A�S�eߟ� ��� $��H���l��i�� =���a�������� ���h�S���'���K� ��o���
��.��R ��v#5o�� ���<�9r �1�U�y� ��8/#/\/��// �/?/�/�/u/�/�/"?�/F?,_>T3 1� I_�/???�?�?�?�/ O�?)O�?&O_O�?�O O�OBO�OfOxO�O�O %__I_�Om__�_,_ �_�_b_�_�_o�_3o �_�_�_,o�oxo�oLo �opo�o�o�o/�oS �ow�6HZ� ����=��a�� ^���2���V�ߏz�� ������]�H���� ��@�ɟd�Ɵ����#� ��G��k���*�d� ů��鯄����1�̯ .�g����&���J�ӿ n�����̿-��Q�� u�ϙ�4ϖ���j��� ��߲�;�������4� �߀߹�T���x��� ��7���[������ >�P�b������!��� E���i��f���:��� ^����������� eP�$�H�l ��+�O�s<Y?k44 1�v?  2l��/2/� V/�S/�/'/�/K/�/ o/�/�/�/�/�/R?=? v??�?5?�?Y?�?�? �?O�?<O�?`O�?O OYO�O�O�OyO_�O &_�O#_\_�O�__�_ ?_�_c_u_�_�_"oo Fo�_joo�o)o�o�o _o�o�o�o0�o�o �o)�u�I�m ���,��P��t� ���3�E�W����ݏ ���:�Տ^���[��� /���S�ܟw� ����� ����Z�E�~����=� Ưa�ï���� ���D� ߯h���'�a�¿�� 濁�
ϥ�.�ɿ+�d� ����#Ϭ�G���k�}� ����*��N���r�� ��1ߓ���g��ߋ�� ��8�������1��}� ��Q���u������4� ��X���|������5 1�M�_��� ;A�_��� ��T�x�% ���j�> �b���!/�E/ �i//�/(/:/L/�/ �/�/?�//?�/S?�/ P?�?$?�?H?�?l?�? �?�?�?�?OO:OsOO �O2O�OVO�O�O�O_ �O9_�O]_�O
__V_ �_�_�_v_�_�_#o�_  oYo�_}oo�o<o�o `oro�o�o
C�o g�&��\� �	��-����&� ��r���F�Ϗj�󏎏 ��)�ďM��q���� 0�B�T����ڟ��� 7�ҟ[���X���,��� P�ٯt����������� W�B�{����:�ÿ^� ������ϸ�A�ܿe�  ��$�^ϿϪ���~� ߢ�+���(�a��υ�� ߩ�D��߳���6 1���zߌ���D�/� h�nߌ�'��K���� ��
���.���R����� �K�������k����� ��N��r� 1�Ugy�� 8�\��}� Q�u��"/�� �/|/g/�/;/�/_/ �/�/�/?�/B?�/f? ?�?%?7?I?�?�?�? O�?,O�?PO�?MO�O !O�OEO�OiO�O�O�O �O�OL_7_p__�_/_ �_S_�_�_�_o�_6o �_Zo�_ooSo�o�o �oso�o�o �oV �oz�9�]o ����@��d�� ��#�����Y��}�� ��*�ŏ׏�#���o� ��C�̟g�🋟�&� ��J��n�	���-�?� Q����ׯ���4�ϯ X��U���)���M�ֿ�q�������7 1� �ߧ����q�\ϕϛ� ��T���x���߮�7� ��[�����,�>�x� �����ߘ�!��E��� B�{���:���^��� ������A�,�e� � ��$���H�����~� ��+��O����H ���h��� K�o
�.� Rdv�/�5/� Y/�}//z/�/N/�/ r/�/�/?�/�/�/? y?d?�?8?�?\?�?�? �?O�??O�?cO�?�O "O4OFO�O�O�O_�O )_�OM_�OJ_�__�_ B_�_f_�_�_�_�_�_ Io4omoo�o,o�oPo �o�o�o�o3�oW �oP���p �����S��w� ���6���Z�l�~��� ��=�؏a����� � ����V�ߟz����'�<��8 1�*�ԟ � �����¯ȟ毁� 
����@�ۯd����� #���G�Y�k����� *�ſN��r��oϨ� C���g��ϋ�߯��� ���n�Yߒ�-߶�Q� ��u�����4���X� ��|��)�;�u����� ������B���?�x� ���7���[������ ����>)b���! �E��{�( �L��E�� �e��/�/H/ �l//�/+/�/O/a/ s/�/?�/2?�/V?�/ z??w?�?K?�?o?�? �?O�?�?�?OvOaO �O5O�OYO�O}O�O_ �O<_�O`_�O�__1_ C_}_�_�_o�_&o�_ Jo�_Go�oo�o?o�o co�o�o�o�o�oF1 j�)�M�� ���0��T�:�L�MASK 1�W��N�����x�XN�O  ������M�OTE  ǌ  ���_CFG ���O�l�PL_�RANG ��q[���A�OWER ��W�y�`�SM_D�RYPRG %�W��%����TA�RT �q���U?ME_PRO������H�_EXEC_�ENB  �t\�GSPD��6�>�;K�TDBY�k��RMz�k�IA_O�PTIONQ���^��INGVE[RS��Ȋ
��o�I_AIRPURO� ��Մ1�m�MT_��Tl��`��OBOT_ISO�LCŌ�-�4�0�^o�NAME����n�OB_CATEGňy�փ̀����سORD_NUM� ?q�*��H769  ��t@�R�d�x�PC_TIMEOUTQ�{ xx�S232��1�ȅj� L�TEACH PENDAN���8����Ƽ ��p�Maintena�nce Cons��r����"���t?No Use��� ��@�R�d�v߈�v���GNPOΐ��8�̥���CH_L����^�J�	���!�UD1:1���R��VAIL!�¥��\��SR  ��ʡ8���R_�INTVAL���\��໮��V_D�ATA_GRP �2�ȅ�� D��PL�/�H�S�>� ȅv���n��������� ��������F4j X�|����� �0TBdf x������/ /*/P/>/t/b/�/�/ �/�/�/�/�/??:? (?^?L?�?p?�?�?�? �?�? O�?$OO4O6O HO~OlO�O�O�O�O�O��O�O __D_́�$�SAF_DO_PULS���p[��OSCAN}���[����SCm�� ��`Xj�W�p�p
���1�`��վQ�r  H��_oo,o>oPo�_�to�o�o�o�o�o����ib2�d�Qy�d�dq�	�T�i @7�FXjtv&y�: ��t�_ @�sTʠ������T D���+�=�O�a�s��� ������͏ߏ����'�9�K��߯�8w�Z�����n�  =��;�o��ʑ��p����
�t��Di_�jaѰ�?X � ���� �U�Q9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ���������	ߗ���2�D� V�h�zߌߞ߰���� �e�� ��$�6�H�Z�@l�~�����}�0�r ��&�������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�� �/�/�/�/�/�/?? +?������ibk?}?�? �?�?�?�?�?�?OO 1O?IROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_��_�_oo&o8o,x� a��Co�o�o�o�o�o �o�o�o"4FX j|���zmo�\��v��+�����	12345�678]2h!B!��%�\1}�k`�T�f�x��� ������ҏ��lo� �1�C�U�g�y����� ����ӟ���	��-� >���a�s��������� ͯ߯���'�9�K� ]�o���@�R���ɿۿ ����#�5�G�Y�k� }Ϗϡϳ����ϖ��� ��1�C�U�g�yߋ� �߯���������	�� -���Q�c�u���� ����������)�;� M�_�q���B������ ����%7I[ m������� �!3EWi{ �������/ ///�S/e/w/�/�/ �/�/�/�/�/??+?@=?O?a?s?�?McE��?�?I/�?�?O�Cz  BpIj_   �H2_b� } �6F
[G�  	�AD�?�O�O�O�O�KDo�<�uO_$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Voho�O�o�o�o�o�o �o�o
.@Rd v�������D#��B�1iA�<�� �iA  �/�I��v,�mA>mAt  6@m�����x`�$SCR�_GRP 1��*P30� �� ��A ��	 Ё�؂�� �1����w��#��J��M�K@G�DC�v���N�G��L�	M-10iA/�8L 12345_67890k@��� 8k@MT20� ͐-C
ș�X��A^H �؁�Z�ǁ'�ǁ�C�G���-�	�v����������ά��H�؀_�܇ǂ���@�5�G���o�A"����������^� �h@,V� � ��B�%@Ɛ������A6@ � � @�@8��N�?��^���H%@q�K��F?@ F�`�£� ���ϲ�������!�� E�0�i����8�h�0ߑߣߵ�B���X� 	���-��Q�<�N�� r���������O� q�3�!�F��]@C��x��B`�8�>����~�6�i�@8���%@���ȗ�'��?�-DA��1a�]�$> �A2�A T{��
i���� (� �  $��H3l)J��Γ���ECLVL  ��A��7�?A���*SYSTE�M*�@V9.10�214 �8/2�1/20�A ��@�z�SER�VENT_T �  $ $S_�NAME !^	 PORT�@!�ROTO! �_�SPD  ���/ TRQ  � 
,#AXISr5!:'2  2c��,#DETAIL_�  l $?DATETI! ERR_COD�#IMP_VEL4@w 	�"TOQ�$�ANGLES�$D�IS��&" G%%�$LIN�" +$R;EC5! ,!O%�i � MRA�! �2 d2IDqX�"�$B  �0�$OVER_L�IMI I �,#O�CCUR5! � �+COUNT�ER!���SF�ZN_CFG5!� 4 $ENA�BL�#ST� "F�LAG"DEBU��3R�!�~3��5!� � 
$MIN�_OVRD�@$�I�� �2�1�5FAsCEe"�1SAF�7MIXEDL�9�!��2ROB%$N�E&APP!��S�HELL�4	� 5$J?@BA�S�#RSR_�5 � $NUM_\y@�  xA1�'�y@2�J3�J4�J5*�J6�J7�J8�'lAgROO � CO��ONLY�$U_SE_AB#xB?ACKENB�  P�IN>0T_CHK�SOP_SEL_��0,Y_PU;Qo1M�_�!OU#PNS@|F PYC�&�0EPM�%�TPFWD_KA�R�! P�!RE$$OPTION�2O$QUE�Y" D�R�YRB$CSTOP�I_AL;SYCEX�+STQ�P�$XTSPM�1i2"MA�1S�TY;TSO
`NBvRDIGQTRI�3\�Q�WINI�M& �8bNRQxf`EN�DNd$KEYSWITCH�S�QZa��THE�PBEAT�M�SPERM_LIE�"�QE� �gU�S�Fd�RS_dDO_�HOM�0ORA/PE�FP !"0�3U ST4�bRC�`OM�#�!�OV_MSJQ ET_IOCMN+Sd�W5a�2ZCHK !�
 D �7qS�U�"�RMP+S� P�O7B$FORCމSWARNk|OM�rP 7�$F'UNC��3U	0}QSAR'`�u2�v3�v}4�q���SC0�O�PL�r�"�XU�NLOeP�$:�E�D� ��SNP�X_AS�2 0·@ADD�0�1$�SIZ�!$VA�R�'MULTIP�RZ��pA�q � $tY[�rC	�B`�"�AC� �ΆFRIF">0S��P�y"t��NF{dODBUS_ADw2��B��&CM�aD�IA�q$DUM�MY15aM�3J�4�J��Sz@  �3 x��"TEqM��8J�SGL��TA>Jp  &�0����@J�����STMT<�Q��PSEGb���BW�P��SHOW���!BAN̐TPSOF�M�9J�0J�~(a�SVC��G�2 ��$PCppP?0-�G3$FB�q-PD�SP�PAFPF��+ VD/��27� ��!A0��@ � ���p���p��	���T���5��6��7��U8��9��A��B��@�p��h ��Ր��F�� �P���T�P���l�P��̩1٩1�1�1� �1�1�1'�1
4�1A�1N��!ǘ�U2��2��2��2̩U2٩2�2�2 �U2�2�2'�24�U2A�2N�3��3��U3��3��3��3̩U3٩3�3�3 �U3�3�3'�34�U3A�3N�4��4��U4��4��4��4̩U4٩4�4�4 �U4�4�4'�44�U4A�4N�5��5��U5��5��5��5̩U5٩5�5�5 �U5�5�5'�54�U5A�5N�6��6��U6��6��6��6̩U6٩6�6�6 �U6�6�6'�64�U6A�6N�7��7��U7��7��7��7̩U7٩7��7�7 �U7�7�7'�74�e7A�7N�L2VP�`=U3" < ƑB
*�� ! x $TOR�QV@�  �"M$ R1 ,L@BQ_W0R��%(T!�p�$S[C�Qp��_U��	 �)�YSL�   � x���7��m��0���`�R�VALAU�5QP�V]�F��ID_L�"%HI�*I�r$FILE1_xSM$BD$s*0��SA21 h�5y E_BLCK��S�"���(D_CPU�)y��)m��3P/b$�p"�`sRR  � PWY0P��6 1LAƑS113�14RUN_FLG(54,14�`/5M14M15HrP4o04� 
�T2�Q_�LI�r  �k@G_Ob�PP�_EDI+Rp�T2 @�3�20�$P�!������TBC2x� �}�8P/0T�Q�1FT'dD5cTDC/0A`a�0@aM	�F.AGTH�"��DDOPGRQH��pERVE(crD5c�rDa��14PG@ �X -$�AL�EN(c�D5c�@`R1A�PF��W_k�#i1�A:$2�GMO�!C�S�DPIZP�F!0Y8�@![DE1U��LACEXrfCC8B���`_MA^�0V8jU@WjQTCVq\�Q@WT�a�Z�U�Zd�/SP]��U@S]�J@`AG��M�T Jjgv�/Ua@U�A2)pp\��5a.SH�JKHfVK@$�ZaU�Zaa�O`J�lra^cJJfcJJncAAL^c�`fc�`�fdm��b5OC�PN1�\P�`�[nP�L
P_��n 2 �1CFb�� `5GROUP ���P�N�0C��~ pREQUIR]B��EBU̓�A�V$T1P2Vq�@@v8�1a��4 \�p�8oAPPRLpCL��
$�0N�xCLO��0�yS:E�y/U�0B]C�� ��0M,@poP�PF��t_MGI��pCx�z �d�lP��BRK�NOLD<��RTMO�1I�$6��uJ�0H�P�dLP fcLPncLP�cLP�cLP%6��7������A>�4� Ir�B�$��U��PATH������H��pr[p�.�SCA�2�L��r�qIN�BUChP�A\�Cf�UMe�	Y�@� `l�&!xA�����������PAYwLOAD�J2LOR_AN$AȓL0�ҙΑޑ�R_F�2LSHRlD�L�OӔ[��i��i�ACRL_�AY�L�U�五gbH��$H��z�FLEX�su �0J�6 P�r@�?
OqO�O �qJ�E  :�O�F@P �#��Oha@P�O�O�LF1#�q����O__0_B_T_��E^_p_�_ �_�_�_�_�_�_�ȩ� �WcHd����o!o3o$"�:jT�Ǌ�Xra Fe���QeZ�3�]ooo �o�`�e�e�e�e�o�o��o�i�2Jt! ���0#5 AT��Hq�PEL�T1p�jOxJ[p VpJE3�gCTRU���TN)�l�@wHAND_V�B��� ׄ" M$��F2�<D��SW !�C�v#� $$M��yM#���2�-�O� �q�K�A@) ���v(!h� �A��#�A1�A@�s��T� #�D1�D@�P �G"0		ST%�2�NC�DY.0�p� T�{����@�#���@��Hg��K�-�G�P�� ������������ʂЂJ�5$ ����� Ʊ�qAS�YM0��Ip0�#wL��P�_n0A�a� t�^�`��~�������ƓJ͜~�ߚ����.��_VI��<(�sM V_UN�2; b#��
�JIez"�z"� ~$4��$�&=��PP�~�_�q�5;�������f�0HR�0�1%��01���2DI@�;sOpO4��10�& ��
��IeA��4�|1�����3��|�0�20 �' � ��M�E���Х2�"�TC0PT����1�`��d����8�1�9T���a $DU�MMY1��$P�S_��RF^�  t�(F�pFLAp�YP2�BB�3$GLB_T�E5]E�0ౡр۰��1( XX�p@wׁST��Vp�SBR�M21_�VRrT$SV_E�R�O��C�CCL�w@�BA�O2,0G�LD EWq) 4\p�1$Y��Z��!WS>`���A�0e�t���AU�E* ��yN P�$GI���}$�A )q��CPq+ Lp\AV�}$F�EIV�NEAR�N��F��Y�TANC�� ? �JOGR�t�� ,^0$JOgINT=�N����C�MSETq-  ">WEvU�:�SA�+1�^Q;�q.� ڥ�U��?�VpLOCK_FO���K0oBGLV��GL:hTEST_XM�pN�QEMP�PRr^buB%`$U��B=�#2*VpS�a+Ob��4*`�a)�ACE�`RS��` $KARP�M>Q3TPDRA�@�d��QVEC4��f�PI�U�a,�aHE,`T�OOLe��cVd�R�E�`IS3�r6�����ACH�P[p-�qO>��3D3���QPSI�r  @�$RAIL_BO�XE=��@ROB�OUd?��AHOW�WAR��tq%@@qROLM0B�u �=t�rp0�bp��ـO_F1��!�@HTML5<D1U� 12�B2qRځ/�^ЀR�`O��a0�R]��Q�p�U;OU�R1 d�@�e�)�v�P�%`$PIPVfN0�rbr2q𫰄a�p�CORD�ED*`6���PXT�V�DQ),0,�O�0 �2 D \@OB��z�*`����C[@����|�SYS��A�DR{�,0�0TCH�:� 3 ,��E�N52��A1a_AT��	����PVWV�A�14 � ��`�BE5PREV_�RT�$EDI}TT�VSHWR1��Fs�� Q< D�0�����$H�EAD�� ����\�KE Q@CPS�PD��JMP��LdD5�0R�g45��T���I_`S{�C���NEp|��TIC)Ke�oM��{A�{HN�A6 @��8��Ñ_GPR�Yvγ�STY	�>qLO�wA ��N� �7 tk 
O�G�%$4��AT=�@Sq�!$@p!=м1HEy0GFPRR�SQU�`X�IB;!�TERC�0����S�8 HP�@.� 0�-���a^�O�0�3F��IZJDAQFE$A�PR��1Ap���.�P9UAဵ_DO�R��XS�PKD6AXI4���s�aURI��@|�{p@�͆��J�_�`߂ET�P3b��5%��F5��AB8D9Hw��UpXR{SR��9l � �M�%�[�8�m�K�[� V�[�d�[�t��Ŗ��� ���Ŷ�����������$!��C6���C�ͯp����qSSC_@� : h�@DS�`��a@SPv0��A	T��L���?��B�ADDRESsB�_�SHIFA�{`_W2CH{�ɁI~@���TU~@I*� �;�RCUSTOT��QVbIj2< �PGh��d�
^j
��qV-����0= \�@�G����o�>�����C���A��~�F��B���TXSCREE���><0��TINA�COP��AT,����? T���@d�߁ �A�@L���ނ��H�[�RRO �Pހ��E��Ŵ��UE�@ ��-��6@S�A߁RS	M?���U��
�D6��00S_S��i�������i�Cb��3� �2?��UEApp2�Bp�GMT� �L�!���@O �_�BBL_BpW�0N�0B ���vOQ�LE�zpE�ތRIGH�BRyD�D�CKGR�0�T����WIDTHHs��ĲUqBAq��UI�pEY�Щ1C6��p�p��bp=l�BACK��0B41�A�0FO�D�LAB��?(�0I<@p#b$UR�qq�YP
�0Hl� D 81�P_����0R P%b/�Hx A�PR�O�0EI��G�� U� �R3b�qL�UM�Ķ�ERVHM��@
P�PF�0�GEu{Q����&��LP4%
�E���)Q'��_(��_(,p^)U5\+6\+7\+8A"���3k��P��F,q�aS��E	US=R�DG <�@�01UERT�ERFOB�ERPRI�mLp�!30�TRIP^qm��UNDOg5H<P`àL0���q����{bްؠ I�� o�G ��T�p�� �&�2OS�1�6R�r�v3�a�AJ�OS^�2Hb�!|aU<!�AK�?��?��<"a�v3OFFTT`�@L�@�3OU@� 1J�@?DgDK�@GUفPfA��C8}ьGSUBb��@N/ SRT�0B�MI���Q�pO�ORBp�ERAUT��DT�I��A9_R��N |]���OWNy0�$S#RC}�����DT`>UR�MPFIy�y��ESP|�G��u#���'rSm�6O� `@WO����=��COP!A$հ{0_YPr�Q.��UWA_�Cra�Q�P�S��Qr;�4��rW� �P?�SHADOW���s"a_UNSC�A�c"c�/cDGD<7q��EGAC�Sd�5��G�Q���'STE���O���t�PE"��VW6Dt�&�RG�6�R �>��jMOVqE}�#A�bANG����f-C�f�3�bLIM_X!Cv'Cv�hq�|��g?06��`"BVqF���CF1VCC��j�S?�C��RA��p�`ϥD��@NFA�Ri@�]�E,�Q>0�G����R:�{0D�E�c�p���p6TG� i�؁ϣ�u��㡹W C% �D#RI�`��aV[�*���S�D�$MY_UBY�$�}�3ϥ~�������Q��P_h8`y���L��BM��$�DEY
�E�Xc ���UMUِX�d����US��˰.0�_R�"B#06��fG�PACIqt�`HQ �dI�-CI��3I����QCRE���1�B�s�I��U ?�PGB�`P�⎐/��sR�0��V�k���B	4�R��R�dSWA�os��@��n�O�!�A(��[�E� U���a��@���sHK��W���aS���Q��c�EANS��P��A�C�sMRCV6X� �- O�pM�C���	��?C����REFb������
r�ِ 0��ꡨ�꡹����A�_;PW�B�o����` ��k�\���x�
b�q3Y ��a��ϒ�1~`�$GROU�� �3��¶�s�pT���х20$ ����0X �V�Ӂ�ֱ���UL��qW�PC%p�X��NT�S+ĔR*� �6��!6���L��_Š��_��k��!�pT�IЙ�Z t@MD>�@AP_HUx��`v��SA�cCMP}�F�����Ų�_��R qty���W�j�X�Ƀr�GF`S[� ��M0����UF�_{�˂��@JʼRO � T�շ����|.��URE9��6�RI;���I&༨�o�o{`FQyFQ'C`wIN�H��xx� V�1,r��A��?�W�|��Q/�0�V큂��LOp'��\ax �����!NSI�IBVIA_�R;�\� �� HDR �)$JO� b�$Z_UP)p>��Z_LOW����@���\(p���P�@�3�9���Ⴐ��'�Q� ���"�]�� 0�PA� �CACH���}�@��퀙�!�P]SC(q%IB�F#���T� ��N|�$HO���� /�%�"f������?�0RQ0!��cPVP��� �H_SIZ�RZ���M��N�Q�MP\r
�qIMG�d��sAD�	�RMRE����WGPM�pND�RP�VASYNBU=F�VVRTD� �W��OLE_2DP,tc�1@C�qUۃ��Q��ECCU{�VEMe�}�d��VIRC��
" {�LA��RQ}0\0֑�AGR�XYZ)��C�W��������A�T�p܂IM��G`��GRABB�1Y�b~� ����^@
�CKLA�S�¡b�Y@_ I 񱵵T��5P@�2��$b��p!�` � ��SP�G�%TQ�RQ�q�P�"x�I�$|���=�BG_LEVE�QL�PKL��"ѥ��GI� NO�Q܁ �a�_HObPRa � �F����E6�S��g]2RO�cA�CCEe@����x4VR�A�y1܂R`� AR�cPA@�>��}D�SREM_BQ$s �p͐JMPU��XAbi$1�$SS(lSFD��S�G�Y@_c  ��S� ���N/D�VLEX�&dbSdqg`��&DR�w$YQqH(`�qH҄�c��P2>h�e� �є`�V��cPMV_PI ��DX�`�@3����I	F&�\rZ�JT�E�@`���H���E�AGAU�?�LOO�d?�JC�BTZ�'B`H +cP�LAN'r��L2��F@w��D?V5Y �WM��~Ppu�T�FS��U �Q�ѥU����V2DbrX�1LRKEZq��1VANC]C`�Rs_O�|`f (�p�8�s$\�3Zr��R�_A3� g 4 ��dovn#p� �݀Sa�ph h��9���.�vOFF�sfW@��,���EA��
� L�SK��MN��q�g� S`��|@c"i �< WJ��=�UM�MYY���n�D6�P�Y!CU��1ѽU�pj $�T�ITV1$PR�8A��OP����SF���Cki �|6���.�BSMO!�l%BXCb�4J�p��ZD�vgm DQx�AL^1#IM; ��0IN�_MSG_Q�S.w ��_p	n%B�w8�%�M� o�XVR"�oI"�pT�5�0ZABC���p��Ƃ��Ӡ
��q%��`VS.� q � w0���=�CTIVeAI�O�b�	s�ITVlLW�DV@
l�"��2� DI�� @�� ��|A��d���N�LSTs���ݰ��7_ST��AA%��DCSCH��r LQp�����~P1��m�W GN����r���_FUN�� �A7ZIP!�s%B� �L8�L|�Ѣ���_ZMPCFʅt�r�9���L�DMY_�LN$pq7�'�˄u $��Q��CMCM��CLCOART_����P�a? $J����D=��¢��u�ǥu����_�����U�X�P�UXEUL ����
�̥
��.�8�>���FTF����k���I�Z�v@_��*�I 7��Y%��D.  w 8 �$R� U�Q��EgIGHe3�x?(�pĚ�0�>p��A$x a�=0�sq�$B������b_SHIYFB�	�RV�PF��&1�	$)0C�ঢ ���d�pl��r�"l���D|ȕ�C �NV:�a	��SPH�0%чy ,�p��ֿ���$S{0DEFA�Un�������������HOT䣐����MIPOWERFL '1�����%�WFD-O�� �� ��Y�~�`1 ���qѾ� L!ip_�EIP5ԑ����j!AF���`�߼�O!FT������f�!��-����.S�!R9MHQp�7�B��f�@o�5�������!OPC3UA�����7�!TPP�@8���yd&���!
PM�p&�pXY����er����J����f��!�RDM-@V��g|
g!R90h2��hV�!
h�~������i��!R�LSYNC &�8�K!ROS̉�r�4:�!
CEL�MT�`��֙k��!	��PSd���l�//!��WASRC6��m�/{/!�USB�|/��nj/�/!S#TMP��/��o�/?@�7?*?`=e�I���KL ?%q� �(%SVCPR#G1`?�:�52�?�?"�03�?�?�04�?�?"�05 O%O�06HOMO"�07pOuO�08�O�O�09�O�K�4~�O �1�?_�1�?=_�1�? e_�1O�_�1:O�_�1 bO�_�1�Oo�1�O-o �1�OUo�1_}o�1+_ �o�1S_�o�1{_�o�1 �_�1�_E�1�_m �1o��1Co��1ko ��1�oe?w2�0~?�0 0�u��1y��������� �Џ	��-�?�*�c� N���r�����ϟ��� ��)��M�8�q�\� ������˯���گ� ��7�"�I�m�X���|� ����ٿĿ�����3� �W�B�{�fϟϊϱ��������k:_DEV� q��M{C:�4���?GRP 2q�����0bx 	�/ 
 ,c��|� <�hߥߌ��߰����� ��#�
�G�Y�@�}�d� ����������d� 1���U�g�N���r��� ��������	��? &cJ����� ����;M4 qX������ /�%//I/0/B// ��/�/�/�/�/�/�/ �/3??W?>?{?�?t? �?�?�?�?�?O�?/O AO�/eOO�O�O�O�O �O�O�O�O_ _=_$_ 6_s_Z_�_~_�_�_�_ �_HO�_'o�_Ko2ooo �oho�o�o�o�o�o�o �o#5Y@}d v�
o����� 1��*�g�N���r��� �����̏	���?� &�c�u����P���ϟ ���ڟ�)��M�4� q�X�j�����˯��� ��%�|��[��� f�������ٿ����� ��3��W�i�Pύ�t��ϘϪ���7�d ���	���	�B�-�f�Qߊߙ�%��߾�>�����у����� ������9�'�]�k� �ߐ���S������� �����;�}�b���+� ��������������C� i�:y�m[� ��� ?�3 �CiW�{�� ��/�///?/ e/S/�/��/�y/�/ �/?�/+??;?a?�/ �?�/Q?�?�?�?�?O �?'Oi?NO`OO9OO �O�O�O�O�O�OAO&_ eO�OY_G_i_k_}_�_ �_�__�_=_�_1oo UoCoeogoyo�o�_�o o�o	�o-Q? a�o�o��o��� ��)��M��t�� =���9���ݏˏ�� %�g�L�����m��� ����ٟǟ��?�$�c� �W�E�{�i������� կ���;�ů/��S� A�w�e���ݯ¿Կ�� ������+��O�=�s� ����ٿc��ϻ����� ��'��Kߍ�r߱�;� �ߓ��߷�������#� e�J���}�k��� �����+�Q�"�a��� U�C�y�g�������� ��'�����+Q? uc�������� �'M;q� ��a����/ /#/I/�p/�9/�/ �/�/�/�/�/?Q/6? H?�/!?�/i?�?�?�? �?�?)?OM?�?AO/O QOSOeO�O�O�OO�O %O�O__=_+_M_O_ a_�_�O�_�O�_�_�_ oo9o'oIo�_�_�o �_oo�o�o�o�o�o 5wo\�o%�!� �����O4�s �g�U���y������� �'��K�Տ?�-�c� Q���u��������#� ����;�)�_�M��� ş����s���o�ݯ� �7�%�[�������K� ����ſǿٿ���3� u�Zϙ�#ύ�{ϱϟ� �������M�2�q��� e�S߉�w߭ߛ߽�� 9�
�I���=�+�a�O� ��s��������� ���9�'�]�K����� ����q��������� 5#Y�����I� �����1s X�!�y��� ��9/0/�	/� Q/�/u/�/�/�//�/ 5/�/)??9?;?M?�? q?�?�/�??�?O�? %OO5O7OIOO�?�O �?oO�O�O�O�O!__ 1_�O�O~_�OW_�_�_ �_�_�_�_o__Do�_ owo	o�o�o�o�o�o �o7o[o�oO=s a�����3 �'��K�9�o�]�� ���̏������#� �G�5�k�������[� }�W�ş�����C� ��j���3��������� ������]�B���� u�c������������ 5��Y��M�;�q�_� �σϥ���!���1��� %��I�7�m�[ߑ��� ���ρ���}���!�� E�3�i�ߐ���Y��� ����������A��� h���1����������� ����[�@�	s a�����! ���9o]� �����/� !/#/5/k/Y/�/��/ �/�/�/?�/?? 1?g?�/�?�/W?�?�? �?�?	O�?Oo?�?fO �??O�O�O�O�O�O�O _GO,_kO�O__�Oo_ �_�_�_�_�__oC_ �_7o%o[oIoko�oo �o�_�oo�o�o3 !WEg��o��o }����/��S� �z���C�e�?���� я���+�m�R���� ��s�������ߟ͟� E�*�i��]�K���o� ������ۯ��A�˯ 5�#�Y�G�}�k���� 	�ڿ������1�� U�C�yϻ���߿i��� e���	���-��Qߓ� x߷�A߫ߙ��߽��� ���)�k�P���� q���������C� (�g���[�I��m��� ����	��� ������ !WE{i���� ���	S Aw���g�� ��///O/�v/ �?/�/�/�/�/�/�/ ?W/}/N?�/'?�?o? �?�?�?�?�?/?OS? �?GO�?WO}OkO�O�O �OO�O+O�O__C_ 1_S_y_g_�_�O�__ �_�_�_o	o?o-oOo uo�_�o�_eo�o�o�o �o;}obt+ M'������ U:�y�m�[�}�� ��Ǐ���-��Q�ۏ E�3�i�W�y�{���ß ��)�����A�/� e�S�u�˟�¯��� �����=�+�a��� ��ǯQ���M�˿�߿ ��9�{�`ϟ�)ϓ� �Ϸϥ��������S� 8�w��k�Yߏ�}߳� ������+��O���C� 1�g�U��y������ ������	�?�-�c��Q�����������$�SERV_MAI�L  �����~��OUTPUT��_��@���RV 2w�  �� (��I���SAVE��TO�P10 2#	 d ���� ��'9K] o������� �/#/5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�?�w�{YPf��FZ�N_CFG w���W~�1GRP 2�7�t ,B   �A'@��D;� B}(@�  B4��RB21VH7ELL�2	w�r�6 7�7�O�K%RSR�O�O�O�O�O _�O3__W_B_T_�_ x_�_�_�_�_�_on?�  ��Ro�Ko]o+bio ���eo�b�`�bg3b2���dultm�bRFHKw 1
`K �o 0YTfx ���������1�,�>�P�LLOMM� `O��QBFT?OV_ENB��+�r�bOW_REG�_UI����IMI_OFWDL�����*E��WAIT�� �i�2����*�wTIM���T��VA��+���_UNcIT����r	LCڀWTRY�r���MON_ALIA�S ?e��2 he���!�3�E�S��� v�������W�Я��� ��ï<�N�`�r��� /�����̿޿𿛿� &�8�J���[πϒϤ� ��a��������"��� F�X�j�|ߎ�9߲��� �����ߥ��0�B�T� ��x������k��� ����,���P�b�t� ����C����������� (:L^	�� ���u� $ 6�Zl~��M ����� /2/D/ V/h//�/�/�/�/�/ /�/
??.?@?�/d? v?�?�?E?�?�?�?�? O�?*O<ONO`OrOO �O�O�O�O�O�O__ &_8_J_�On_�_�_�_ O_�_�_�_�_o�_4o FoXojo|o'o�o�o�o �o�o�o0B�o Sx���Y�� ����>�P�b�t� ��1�����Ώ��򏝏 �(�:�L���p����� ����c�ܟ� ��$��Γ�$SMON_�DEFPROG �&���N�� &*S?YSTEM*+�o�����?=�R�ECALL ?}�N� ( �}!�xyzrate �124=>169�.254.��12�0:14636 ���ĥ�����}
��1 ��ǯٯj�|� ��!���;�M�_����� }:copy� frs:ord�erfil.da�t virt:\�tmpback\`���qσϕ�}1*�mdb:*.*?πQ�ʰ]��� ��%�5x*�:\��4���ǲ���q߃ߕ�}6*�a 2�D�·a�����)� ;�����p����B� ��]��� ��%߸��� [�l�~�����4�F���P����!��� �������k}�����19ȱL^�&�����m�$�m�d:picksi�m_part1.;tp��emp��F ��/��?���o/�/�/&tpdisc 0N/GI/�[/�/�/?#tpconn 0 �/ �/�/h?z?�?1Q?@G?Y?�?�?O�52�omay��?ڳ�?qO�O�O(K27OIO[O�O�O_�Ld3O�O�O h_z_�__1R�OH_Z_ �_�_o"/4/F�_�_ oo�o�o&8oJo\o�o �o$o�o�o�ok} ��o�oFX���  2��g�y���� �B�T����	��.� ��ҏ�u����,�>� 7�b������ş>� ݟn�����%�8E�G `��������˯^ o���������A�\�� ���$���ѿZ�k�}� �Ϣ�3�G�د�����  �2���V�g�yߋߞ� ��9�Կ����	��.����R��u����$�SNPX_ASG 2�������  �0�%�����  �?���PARAM� ���� W�	��P��9��1������OFT_KB_CFG  �����OPIN_SIMW  ��,����������RVNO�RDY_DO  �6�b���QST_P_DSBv�,�|��SR �� � &0�Q���G�TOP_ON_ERR����|�PTN ��ޯ �A�RI?NG_PRM����VCNT_GP �2x�.���x 	 
	��0T���VD� RP 1�/�E��7�� �����//1/ C/U/g/y/�/�/�/�/ �/�/�/	??-???Q? c?�?�?�?�?�?�?�? �?OO)OPOMO_OqO �O�O�O�O�O�O�O_ _%_7_I_[_m__�_ �_�_�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/A hew����� ���.�+�=�O�a� s���������͏�� ��'�9�K�]�o��� ������ɟ۟���� #�5�G�Y���}����� ��ůׯ�����F� C�U�g�y��������� ӿ��	��-�?�Q��c�mPRG_CO7UNTW����'ENB���M��Y����_UPD 1>4T  
xϣ� ��/�X�S�e�wߠ� �߭߿��������0� +�=�O�x�s����� ���������'�P� K�]�o����������� ������(#5Gp k}�����  �HCUg� ������� / /-/?/h/c/u/�/�/ �/�/�/�/�/??@? ;?M?_?�?�?�?�?�? �?�?�?OO%O7O`O�[OmOO�O�O�O��_INFO 1�����P	 ��O__@_+Y@�l�@I�l?�Z�F_-S�̵���5Au��9	�]�Ǝ��@�K]A����@CP A!"� ?�nn_�A �D5Oy����C���(�$6�T5+����Q� 8��h�Ca��.�~:��1５����YSDEBSUG������@d���
`SP_PASS��B?kLOG� �F�  ��@�X�O  �����AUD1:�\Hd�NIb_MPC Nm���o�o���a�o� ���fSAV �Qi��2Qqa�b�E��hSV�kTEM�_TIME 1�Qg� 0�����Ļ�h2_�A[vME?MBK  �����q`qo�� �X;|��� @ ��C�"�G�W��z���Y��a �{@}q ��я�����+�=�O�a�s��D�{����� ß՟�����/�i�e>�c�u��������� ϯ����)�;�M��_�q���������\uSK�p�x�������V�1�@|��2,�6W�AW΀ Tý�hi��Ϧ�(��!�������� ����-�g  �-���0�� s߅ߗߋ�Xπ���� ����(��@$,�P� D�t��������� ����(�:�L�^�p��������������T1�SVGUNSPD�2e 'e���2�MODE_LIMC �vvq b��2���Qm��ASK_OPTION`t�y aS_DI+`?ENB  b�e�sBC2_GRP 2ܵc|r�[R��C�����BCC�FG �7| q(��` M_VAf�w�� ����///R/ =/v/a/�/�/�/�/�/ �/�/??<?'?`?K? �?�?8Ձ<�?�?�?�? p?�?+OOOO:OsO~ �O�th@�O�O�O�O�O 	_�O-__=_?_Q_�_ u_�_�_�_�_�_�_o )ooMo;oqo_o�o�o �o�o�o�o�h�0 3EW�o{i�� �������A� /�e�S�u�w������� �я���+��;�a� O���s�����͟��ݟ ߟ�'��K�c�u� ������5�ۯɯ�� ��5�G�Y�'�}�k��� ��ſ��տ׿��� C�1�g�Uϋ�yϛ��� ������	���-��=� ?�Q߇�u߫�a����� �����;�)�K�q� _���������� ��%��5�7�I��m� ��������������! E3iW�{� ������#5 Sew����� ��//�=/+/a/ O/�/s/�/�/�/�/�/ ?�/'??K?9?[?�? o?�?�?�?�?�?�?�? �?OGO5OkO!�O�O �O�O�OUO�O�O_1_ _U_g_y_G_�_�_�_ �_�_�_�_�_	o?o-o coQo�ouo�o�o�o�o �o�o)M;] _q����O�� �%�7��[�I�k��� ���Ǐُ�����!� �E�3�U�W�i����� ß���՟����A� /�e�S���w������� ��ѯ���+��C�U� s����������˿��߿���3��$TB�CSG_GRP �2����  �3� 
 ?�  ^�p�Z� ��~ϸϢϴ�������$�7�>�E�d�0 �S�?3�	 _HCA�"�>l�~"�CS�BpV���ߙ�c�u߇���B��$�>�����"�B�l����)�A����c��G�"�;�B�)�+�Q�G��_��A3�"�Q���T��Ѩ��@�����'�:�� �e���M�_��������?�ff�� ��	�V3.00V�	Omt2 * @2�$��<3�GƯ� [ -\  aq��7�J2>��E���CFG� !��O� �R��
���0�0Vd �d�u���� ��///P/;/t/ _/�/�/�/�/�/�/�/ ??:?%?^?I?�?m? ?�?�?�?�? OOV� p�O/OAO�?tO_O�O �O�O�O�O�O�O_(_ :_L__p_[_�__�_ �_3���_���_oo Io7omo[o�oo�o�o �o�o�o�o3!W Egi{���� ����-�S�A�w� e�����m�ŏ׏���� ��=�+�a�O���s� ����͟ߟ����� 9�'�]�o�����M��� ��ۯɯ����5�#� Y�G�}�k�������׿ ſ�����C�1�S� U�gϝϋ��ϯ����� 	����?��W�i�{� %߫ߙ߻߽������ )��M�_�q��A�� ���������%��� 5�[�I��m������� ��������!E3 iW�{���� ��/?AS �w������� /��O/=/s/a/�/ �/�/�/�/�/??�/ %?K?9?o?]?�?�?�? �?�?�?�?O�?!OGO 5OkOYO�O}O�O�O�O �O�O_�O1__U_C_ y_g_�_�_�_�_�_�_ �_o	o+o-o?ouo� �o�o�o[o�o�o�o ;)_M��� �w�����7� I�[��'�������� ُǏ����3�!�W� E�{�i���������ß �����A�/�e�S� u����������ѯ� ��o1�C��o����s� ����Ϳ��ݿ��'� 9�K�	�ρ�oϥϓ� �������Ϲ�#��3� 5�G�}�kߡߏ��߳� ��������C�1�g� U��y�������� 	���-��Q�?�a��� u���%�W��������� M;q_�� �����# %7m��]� ���/�/!/3/ i/W/�/{/�/�/�/�/ �/?�//??S?A?w? e?�?�?�?�?�?�?�? OO=OOO��gOyO�O 5O�O�O�O�O�O�O_ 9_'_]_o_�_�_Q_�_�_�_�_�_�^  %`)c )f=o)b��$TBJOP_�GRP 2"�U��  K?�)f	Ub\c$cl���P���pJ�`�xe � � � � ���`�)d @�%`tb	 �CA����f��SC��q_)eta�b333�f��oz=�_�C?S�?���1ru`B�;pp�gLWw�o��o?�a�u��z<;؄-r����u=��)eB��wC�  D�a�o#�-�?;��Bl�`2uǦff�n�)eA�䇇�w��>���ͭ�����;ǎ���@fff��b�x]���A����p����9�ˌ�X��@�o�폎�����%�x�ɟۛ;�����@�o���{���� 9�1�g�Y�C�Q���� ��E�ϯ�ӯ��@� �կ_�y�c�q���п�ct�)f��	�V3.00zcmt2��*�yd$a�)�4� F�� G9| G�v��G�/�G��� H�@H,��H.��HC�� HYA@Hn���H�� H��� H�Y@H��`H���H�c��H��H̿��H�nD�G� G.A GKm� Gh� G����G�x�G���G���G�:��G�ЀG�f��G���G���\��H
_�H���H��H� @�H'�d����=L��=#�!
������)b3o�j+�)f/�?�߀�f�d�RcESTPA�RS�hn`RcHR���ABLE 1%*ci�)d_�D�Q �@$�_�_�_ب(g0a_�	_�
_��_ؾ�)a_�_�8_�����RDI��ma�����������O�������������S��kc I���� ������*<N `r������ �Hm����lb��C ,�>�P�b�� �2�D��V�h��)NUM [ �Uma�`�1` �����_CFG &+��a�@U`IMEBF_�TT�Ѻkc��T&V�ER�Uj&T#R� 1'�� 8$&�)b$`�! �PN  �/�/�/�/�/	? ?-???Q?c?u?�?�? �?�?�?�?�?<OO)O rOMO_OuO�O�O�O�O �O�O�O__%_7_I_ [_m__�_�_�_�_�_ �_4oo!ojoEoWomo�{o�o�o�o�oҗ!_�!�&@�%��MI__CHAN`' �%� .sDBGLVL�`'�%��1pETHERAD ?���p�/��o�o�x�y�1pROUT~ !�!�t��|?SNMASKyx�#>�q255.?���=�O�a�Á�OOL�OFS_DI����ecyORQCTRL (�+��0�ߍTΏ��'�9�K�]� o���������ɟ۟� ���#�3�͏V�E�z��~�PE_DETA�IWx��PGL_C�ONFIG .�)"!��/ce�ll/$CID$/grp1~�����*�<����g�y� ��������P����	� �-�?�οc�uχϙ� �Ͻ�L�^�����)� ;�M���q߃ߕߧ߹� ��Z�����%�7�I� ������������M}n��!�3�E�W� i��k���p��m��� ������ g�DV hz��-��� �
.�Rdv ���;���/ /*/�N/`/r/�/�/ �/�/I/�/�/??&? 8?�/\?n?�?�?�?�? E?�?�?�?O"O4OFO �?jO|O�O�O�O�OSO �O�O__0_B_�Of_�x_�_�_�_�_�_͠��User V�iew �}}1�234567890oo'o9oKo]oedX�`£�o���Y2�Y b_�o�o�o�o!�o�o�R3�oo��� ��(��n4^#� 5�G�Y�k�}�����n5�׏�����1���R��n6Ə������@��ӟ�D���n7z� ?�Q�c�u����������n8.����)�;��M���n�t� l�Camera �Z꯳�ſ׿������E��7�I�[�ou���ϙϫϽ���ŉ   ���i���1�C�U�g� y� ϝ߯�������� 	��-�?�f����]y �ߋ���������� 	��-�x�Q�c�u��� ����R�d��B���	 -?Q��u�� �������� d��˰ew��� �f��/R+/=/ O/a/s/�/,��y�/ �/�/�/??)?�M? _?q?�/�?�?�?�?�? �?�/d�-��?;OMO_O qO�O�O<?�O�O�O(O __%_7_I_[_Od� ��O�_�_�_�_�_o �O%o7oIo�_moo�o �o�o�on_�W9So ,>Pb	os� �Qo�����(�:�ɪ	��0�u��� ������Ϗv��� �;�M�_�q�����<� N�����9�� ��$� 6�H��l�~���۟�� Ưد��������� ��Z�l�~�������[� ؿ���G� �2�D�V� h�z�!�[�n������ ����� �ǿD�V�h� �όߞ߰������ߍ� ����}�2�D�V�h�z� ��3߰��������
� �.�@�R��ߟ�F�� �������������� .@��dv��� �e��Ų+U
. @Rd��������//*/�  �	Y/k/}/�/ �/�/�/�/�/�/?;   //7/U?g? y?�?�?�?�?�?�?�? 	OO-O?OQOcOuO�O �O�O�O�O�O�O__ )_;_M___q_�_�_�_ �_�_�_�_oo%o7o�Io[omoo�o#<  }
� (  �M ( 	 �o�o�o �o�oC1SU�g������j?: �y*�<�N� �r���������̏� �����a�>�P�b� t�����ߏ��Ο��'� ��(�:�L�^����� �����ʯܯ� �� $�k�}�Z�l�~�ů�� ��ƿؿ���C� �2� Dϋ�h�zόϞϰ��� 	�����
�Q�.�@�R� d�v߈����Ͼ����� )���*�<�N�`�� ������������� �&�m�J�\�n���� ����������3�E�" 4F��j|��� ���S0B Tfx����� �//,/>/P/� ��/�/�/��/�/�/ ??(?o/L?^?p?�/ �?�?�?�?�?�?5?O $O6O}?ZOlO~O�O�O8�O�?�p@ �B�O��O_�C�G�`���#frh:\tp�gl\robots\m10iaAS_8l.xml�O e_w_�_�_�_�_�_�_�_on��o>oPo boto�o�o�o�o�o�o �oo:L^p ������� � �6�H�Z�l�~��� ����Ə؏����� 2�D�V�h�z������� ԟ����	�.�@� R�d�v���������Я �����*�<�N�`� r���������̿޿� ��&�8�J�\�nπ� �Ϥ϶��������� X�VA �O+P<�< )P ?� ��A���9�[߉�oߑ� �ߥ����������=� #�E�s�Y�����������6�$TP�GL_OUTPU�T 1	A	A !�-�B�T� f�x������������� ��,>Pbt ������-�!�����2345678901); M_g�2��� �����/0/B/T/f/�}p/�/�/�/ �/�/x/�/?(?:?L? ^?p??~?�?�?�?�? �?�?�?$O6OHOZOlO OO�O�O�O�O�O�O �O
_2_D_V_h_z__ �_�_�_�_�_�_�_�_ .o@oRodovo�o o�o �o�o�o�o�o< N`r�.�� �����"�J�\� n�����*���ȏڏ�������}�F�X� j�|�������@#�՟��)� ( 	 ��
�@�.�d�R� ��v��������Я� ��*��N�<�^���r� ����̿���޿ �� �J�8�n����8� vϨϺ͒�������� $��
��U�g��sߝ� w߉�����C����� �Q�c�=����߁� ��i������;�M� ��5�����/������� ��_�q�7I��Q Yk��%�� ��3i{� ��K����/ //�/e/w//�/�/ �/�/�/A/�/?+?�/ O?a?;?M?�?�/?�? �?y?�?O�?OKO]O �?aO�O-OO�O�O�O �O_oO�OG_�O3_}_ �_i_�_�_#_�_�_o �_1oCooOoyo�_�_ �o�o[o�o�o�o�o- ?�ocua�������)WG?L1.XML��(���$TPOFF_�LIM ��������6�N_S]V>�  ��P��P_MON 2���R�����2�2�STRTCHK' 3��P�C�9��VTCOMPAT�e��T�VWVAR� 4���i� KƏ *�I����:�_DEFPR�OG %��%�MAIN  T�Ld�T1A�3�_D?ISPLAYE����Z�INST_MSwK  �� ��?INUSER叜��LCK�QUI�CKME{��Z�S7CRE1�����?tpsc����L�Q�P�b�_f�ST��P�RACE_C_FG 5���uI�	3�
?���?HNL 26i�b�ѡ� ?���)�;��M�_�q�������IT�EM 27� ��%$12345�67890ؿ� � =<���"� G !(�0�<�� u�3�ֿ��������0� ��T�f�/ߊ�J߮�Z� �������4�>߸� b��4�F��j����� ��l��������^�� ����*�x������ ���6�H�l�,�� Pb��x��<�  �D�(�4� ��N����@  /dv�/$/�~/ �/��//*/�/N/? r/2?D?�/Z?�/�/�? ?�?&?�?�?~?n?�? �?�?�?0O�?�O�O�O "O�OFOXOjO�O�O:_ `_r_�O~_�O__�_ �_T_o&o�_2o�_�_ �o�_�oo�o�o>o�o bo�o=�oX�oh� ��(:L�p �B�T��x��� � ����6����l���� ��k�Ə��ꏪ��� ��ҟD�V����S��8|��$��  ���$� ɡ{�r�
 �������үS�UoD1:\߬��6��R_GRP 19�Ż� 	 @{�*�<�&�\�J���n��������˿ٺ���߯��'��?�  B�T�>�t�bϘφ� �Ϫ���������:߀(�^�L߂�pߒ߸�	������4�SCBw 2:@� -� *�<�N�`�r�������*�UTORIAL ;@�Ư�/��V_CONFIG <@�ġx�¯d���OUTPUT �=@�U��� p�����������  2DVhz�R�� ����� 2 DVhz���� ���
//./@/R/ d/v/�/��/�/�/�/ �/??*?<?N?`?r? �?�?�/�?�?�?�?O O&O8OJO\OnO�O�O �?�O�O�O�O�O_"_ 4_F_X_j_|_�_�O�_ �_�_�_�_oo0oBo Tofoxo�o�o�_�o�o �o�o,>Pb t���o���� ��(�:�L�^�p��� �����ʏ܏� �� $�6�H�Z�l�~����� >�P��������(� :�L�^�p��������� ��ܯ� ��$�6�H� Z�l�~�������ůؿ ���� �2�D�V�h� zόϞϰ���ӿ���� 
��.�@�R�d�v߈� �߬߾��������� *�<�N�`�r���� ����������&�8� J�\�n����������� ������"4FX j|������� �0BTfx �������/ /,/>/P/b/t/�/�/ �/�/�/��/??(? :?L?^?p?�?�?�?�?|�?������? �?�1�?&OɟJO\OnO �O�O�O�O�O�O�O�O _"_�/F_X_j_|_�_ �_�_�_�_�_�_oo 0oA_Tofoxo�o�o�o �o�o�o�o,=o Pbt����� ����(�9L�^� p���������ʏ܏�  ��$�6�G�Z�l�~� ������Ɵ؟����  �2�C�V�h�z����� ��¯ԯ���
��.� ?�R�d�v��������� п�����*�<�M� `�rτϖϨϺ����� ����&�8�I�\�n� �ߒߤ߶�����������"�4�C��$TX�_SCREEN �1>�5�0�}�C����������u�2Ft�!� 3�E�W�i�{������ ����������/�� Sew���$� H�+=O� �������V /z'/9/K/]/o/�/ ��//�/�/�/�/? #?�/�/Y?k?}?�?�? �?*?�?N?�?OO1O�COUO�?yO�$UA�LRM_MSG k?c��p� qO FګO�O�O�O__6_ )_;_Y___�_�_�_�_��_�ESEV  �M
f�BECFoG @c�m��  F�@�  }A:a   B�F�
 �_M�c�moo �o�o�o�o�o�o�o�!/waGRP 2�A k 0F�	 �Woy�@I_BB�L_NOTE �B jT��#lM�h�O�,`�r�DEFPRO�@%��K (%MAINz�}%�_�� ?�*�c�N���r�����ਏ�̏��{FKE�YDATA 1C<c�cpp /gF�fi�{�R��������,(���F�ҐOI�NT ER��?DIRECTB`4���IN,�D�F�[CHOICE]p�~�[LIST�� Ư��ܯ�կ���6� H�/�l�S�������ƿ����ѿ�� ϋ����/frh/gu�i/whitehome.png)��g�yϋϝϯπ  >A�pointR��Ϡ����+ߺ�@�direc��g�yߋ�h�߯ߺ�@�inQ߀������0�;�E�choicQ�o��������@�lis ��a���	��-�?���arwrg��w��� ������N�����  $6H��l~�� ��U�� 2 D�hz���� �c�
//./@/R/ �v/�/�/�/�/�/_/ �/??*?<?N?`?7� e?�?�?�?�?�?�?�/ 
OO.O@OROdO�?�O �O�O�O�O�OqO�O_ *_<_N_`_r__�_�_ �_�_�_�__o&o8o Jo\ono�_�o�o�o�o �o�o�o�o"4FX j|����� ���0�B�T�f�x� �������ҏ���� ��,�>�P�b�t���� ����Ο��������:�L�^�p�����/�����:����ʯܯ�Ư�"���,�S��w�^����� ��ѿ������+�� O�a�Hυ�lϩϻϢ� �������'�9� �]� D߁ߓ�r?�������� ��� �5�G�Y�k�}� ���0���������� ���C�U�g�y����� ,���������	- ��Qcu���: ���)�M _q����H� �//%/7/�[/m/ /�/�/�/D/�/�/�/ ?!?3?E?�/i?{?�? �?�?�?R?�?�?OO /OAO�?eOwO�O�O�O �O�O���O__+_=_ O_VOs_�_�_�_�_�_ �_n_oo'o9oKo]o �_�o�o�o�o�o�ojo �o#5GYk�o ������x� �1�C�U�g������ ����ӏ������-� ?�Q�c�u�������� ϟ�󟂟�)�;�M� _�q��������˯ݯ ����%�7�I�[�m� ������ǿٿ������@���@���:�L�^�6��ϒ�l�,~���v��� �����A�(�e�w� ^ߛ߂߿��߸����� �+��O�6�s�Z�� ����������O'� 9�K�]�o��������� ����������5G Yk}���� ���1CUg y��,���� 	//�?/Q/c/u/�/ �/(/�/�/�/�/?? )?�/M?_?q?�?�?�? 6?�?�?�?OO%O�? IO[OmOO�O�O�ODO �O�O�O_!_3_�OW_ i_{_�_�_�_@_�_�_ �_oo/oAo�eowo �o�o�o�o�_�o�o +=O�os�� ���\���'� 9�K��o��������� ɏۏj����#�5�G� Y��}�������şן f�����1�C�U�g� ����������ӯ�t� 	��-�?�Q�c�򯇿 ������Ͽ�󿂿� )�;�M�_�q� ϕϧ� ��������~��%�7ߠI�[�m��V`��}�V`�����@���ݦ������,�� 3���W�>�{��t�� �����������/�A� (�e�L����������� ���� =$a sRo������  �'9K]o� ������� #/5/G/Y/k/}//�/ �/�/�/�/�/?�/1? C?U?g?y?�??�?�? �?�?�?	O�?-O?OQO cOuO�O�O(O�O�O�O �O__�O;_M___q_ �_�_$_�_�_�_�_o o%o�_Io[omoo�o �o2o�o�o�o�o! �oEWi{��� ������/�6 S�e�w���������N� �����+�=�̏a� s���������J�ߟ� ��'�9�K�ڟo��� ������ɯX����� #�5�G�֯k�}����� ��ſ׿f�����1� C�U��yϋϝϯ��� ��b���	��-�?�Q� c��χߙ߽߫����� p���)�;�M�_��� ������������p�����p����,�>��`�r�L�,^��V������ ����!EW>{ b������ �/S:w�p �����//+/ =/O/a/p�/�/�/�/ �/�/�/�/?'?9?K? ]?o?�/�?�?�?�?�? �?|?O#O5OGOYOkO }OO�O�O�O�O�O�O �O_1_C_U_g_y__ �_�_�_�_�_�_	o�_ -o?oQocouo�oo�o �o�o�o�o�o); M_q��$�� �����7�I�[� m���� ���Ǐُ� ���!��E�W�i�{� ������ß՟���� �/���S�e�w����� ��<�ѯ�����+� ��O�a�s��������� J�߿���'�9�ȿ ]�oρϓϥϷ�F��� �����#�5�G���k� }ߏߡ߳���T����� ��1�C���g�y�� �������b���	�� -�?�Q���u������� ����^���);hM_6�a�6�����������,�� 7[mT�x� ����/!//E/ ,/i/{/b/�/�/�/�/ �/�/�/??A?S?2� w?�?�?�?�?�?���? OO+O=OOOaO�?�O �O�O�O�O�OnO__ '_9_K_]_�O�_�_�_ �_�_�_�_|_o#o5o GoYoko�_�o�o�o�o �o�oxo1CU gy����� ���-�?�Q�c�u� �������Ϗ��� ��)�;�M�_�q���� ����˟ݟ����%� 7�I�[�m����h?�� ǯٯ�����3�E� W�i�{�����.�ÿտ ����Ϭ�A�S�e� wωϛ�*Ͽ������� ��+ߺ�O�a�s߅� �ߩ�8��������� '��K�]�o���� ��F��������#�5� ��Y�k�}�������B� ������1C�� gy����P� �	-?�cu@�����������������/-�@/R/,&, >?�/6?�/�/�/�/�/ ?�/%?7??[?B?? �?x?�?�?�?�?�?O �?3OOWOiOPO�OtO �O�O���O�O__/_ A_Pe_w_�_�_�_�_ �_`_�_oo+o=oOo �_so�o�o�o�o�o\o �o'9K]�o ������j� �#�5�G�Y��}��� ����ŏ׏�x��� 1�C�U�g��������� ��ӟ�t�	��-�?� Q�c�u��������ϯ �󯂯�)�;�M�_� q� �������˿ݿ� ��O%�7�I�[�m�� ���ϵ���������� ��3�E�W�i�{ߍ�� ������������/� A�S�e�w���*�� ����������=�O� a�s�����&������� ��'��K]o ���4���� #�GYk}� ��B���// 1/�U/g/y/�/�/�/ >/�/�/�/	??-???��A;�����j?|?�=f?�?�?�6,�O�?�OO�? ;OMO4OqOXO�O�O�O �O�O�O_�O%__I_ [_B__f_�_�_�_�_ �_�_�_!o3o�Woio {o�o�o�o�/�o�o�o /A�oew� ���N���� +�=��a�s������� ��͏\����'�9� K�ڏo���������ɟ X�����#�5�G�Y� �}�������ůׯf� ����1�C�U��y� ��������ӿ�t�	� �-�?�Q�c��ϙ� �Ͻ�����p���)� ;�M�_�q�Ho�ߧ߹� ���������%�7�I� [�m��������� �����!�3�E�W�i� {�
������������� ��/ASew� ������ +=Oas��& ����//�9/ K/]/o/�/�/"/�/�/ �/�/�/?#?�/G?Y? k?}?�?�?0?�?�?�? �?OO�?COUOgOyOЋO�O�O���K�>������O�O �M�O _2_V,oc_ o�_n_�_�_�_�_�_ oo�_;o"o_oqoXo �o|o�o�o�o�o�o �o7I0mT�� �������!�0O E�W�i�{�������@� Տ�����/���S� e�w�������<�џ� ����+�=�̟a�s� ��������J�߯�� �'�9�ȯ]�o����� ����ɿX�����#� 5�G�ֿk�}Ϗϡϳ� ��T�������1�C� U���yߋߝ߯����� b���	��-�?�Q��� u��������� ��)�;�M�_�f�� ������������~� %7I[m���� ����z!3 EWi{
��� ����///A/S/ e/w//�/�/�/�/�/ �/?�/+?=?O?a?s? �??�?�?�?�?�?O �?'O9OKO]OoO�O�O "O�O�O�O�O�O_�O 5_G_Y_k_}_�__�_��_�_�_�_oo�$�UI_INUSE�R  ����@a� �  o$o_MENHIST 1D@e�  �( M`��(/�SOFTPART�/GENLINK�?current�=menupage,153,1_o0�o�o�o�'�o�n71�oSew��Qy)�eedit�bMAINB���p��,�`422��]�o�����4�e,�2�oޏ�����R� �>�P�b�t�����'� ��Ο�������:�@L�^�p��������4� �a4�ѯ�����+� .�O�a�s�������8� Ϳ߿���'϶�ȿ ]�oρϓϥϷ�F��� �����#�5���Y�k� }ߏߡ߳�B�T����� ��1�C���g�y�� ����אָ����	�� -�?�Q�T�u������� ����^���); M_������� �l%7I[ ������� z/!/3/E/W/i/� �/�/�/�/�/�/���� ?/?A?S?e?w?z/�? �?�?�?�?�?�?O+O =OOOaOsO�OO�O�O �O�O�O_�O'_9_K_ ]_o_�__�_�_�_�_ �_�_o�_5oGoYoko }o�oo�o�o�o�o�o �/
?CUgy� ��o����	�� ��Q�c�u������� :�Ϗ����)��� M�_�q�������6�H� ݟ���%�7�Ɵ[� m��������D�ٯ�����!�3���$�UI_PANED�ATA 1F����i� � 	�}c/f�rh/cgtp/�flexdev.�stm?_wid�th=0&_height=10�����ice=TP&�_lines=3���columns�=4��fon��4�&_page=d�oub��1E�!v)�prim��  }�8�J�\�nπ��� )�ϸϟ�����  ����6��Z�l�S߀��wߴ��߭���!v���     �v"��>/FRH/VI�SION/VRF�RMN.STM?�_imӰonly�=1ǰilter�shown��A�eOd=1 ��̿2���dual���$� ��������/���S� :�w���p��������� ����+OaH����k����� �%xI��m ����.�� �!//E/W/>/{/b/ �/�/�/�/�/�/�/?/?� �4?l?~?�? �?�?�??�?]O O 2ODOVOhO�?�O�O�O �O�O�O�O�O__@_ '_d_v_]_�_�_�_�_ C?U?oo*o<oNo`o �_�o�?�o�o�o�o�o io8\C� �y������ �4�F�-�j��_�_�� ��ď֏���M��0� �oT�f�x�������� ҟ������,��P� b�I���m�������� ǯ�w����L�^�p� ��������ʿ=�� � �$�6�Hϯ�l�~�e� �ω��ϭ������� � �D�V�=�z�aߞ߰� #�5�����
��.�@� ��d�׿������� ��I������<�#�`� r�Y���}������������&J������T������) {��8J\n �������� /�4//X/j/Q/�/ u/�/�/�/�/x�������$UI_POSTYPE  ���� 	 ��/K?2QUICKMEN  );�8?N?0REST�ORE 1G���  �	�/���?�3�?��m�?O+O=OOOaOO �O�O�O�O�OpO�O_ _'_9_�?F_X_j_�O �_�_�_�_�_�_o#o 5oGoYokoo�o�o�o �o�o�_�o�ozoC Ugy�.��� ����-�?�Q�c� ���������� ��)�̏M�_�q��� ��8���˟ݟ���� � �2���m������ ��X�ٯ����!�3��֯W�i�{�����Y7S�CREi0?n=�u1sc�0�u2ڴ3ڴ4ڴ5*ڴ6ڴ7ڴ8ڱ��wTAT%=� }3<��:USER�����Ӵksܳm�3m�4�m�5m�6m�7m�8�m�0NDO_CFG H);d c0�PD�W���None\2N�_INFO 1I��5�{00%��� x�
�K�.�o߁�dߥ� �ߚ��߾������5��G�*�k�R<��OFF?SET L)9�x�@��0H������� ����(�U�L�^��� b������������� $6��~?�p��
����UFRA_ME  @������RTOL_AB�RT���ENB� GRP 1M��9z1Cz  A�ec��cu��@����h0U/���MSK  h2�N�%����%Rs/ _EV�N2$�ƈ&��2�N��
 h���UEV!td�:\event_�user\w/� C�7�/�B�F<�!S�P�!�'spot�weld=!CA6????�0b$!b/ �/�?�?�7!�?�?�? OAO�?�?wO"O�OFO XOjO�O�O_�O�O�O O_>_s__0_f_�_�_ �_�_�_o�_9oKo�_�o�o,o�oPobj�&W�RK 2OXɶ8�o	 �o@R -v�c���� ���*��N�`�;� ����q���̏��ݏ����$VARS__CONFI��P�� FP@���C7CRG��S��Z�@�9�D�B�BeH�p����C����їϑ?��U�M�RK2Y���)B�	��C�X�1�: SC130E�F2 *3�7�@�����ch �5B�l���A@��CȐ�' �����9����ȯ���������ӑ��	�Z���? B���u��� z����᯾����Ϳ ��*��'�`Ϸ�A� �ρϓ�������X�TCCc�ZR�4�h�pa��'�GF,���![�� �a 2�34567890�1q�y�'9�n��� n߰ߘ#����j������B��Ӗ ��ϑ:�o=L{��!p�  �p��ia/[�ߤԆ� ����������)�;� (�:�q��p����� ������%�I�[� H���{��������|"�S�SELEC�$�!?�AVIA_[WO�`\T)_>ff,		�= �>;G�P �R'	��RTSYNCS�E�j��n�eWINURL ?u��R����� //"�ISION�TMOU�/ ��*%c�]S۳�S�۵@/� F�R:\,#\DAT�As?MЄ� M�Ck&LOGx/  � UD1k&EX��/��' B@� ���"�!D�ESKTOP-M?C6FJ6K�/�#�?%?�le � �n6  ���x�f�"�� -�N5�K�   =�C��w1��t0� �(TRAIN�/H҆2��bd�3pw5{4� #`�"'(��^]� (���9M�� OO+O=OOO�OsO�O �O�O�O�O�O�O_$(STAT _'�@ �z�b_t_�_�h$�_\�_'%_GES#`]�;��0 �
��|�R�WHOMINV _aS۾�`�b"(���C�ז&�W�JMPERR 2=b]�
  =�j ho^l��o�o�o�o�o �o�o.<m`lr�S_� REV �cO^#�LEX�Td�7��1-e�_VM�PHASE  �j���&�OFF�o_ENB  �\�	P2R$eS�K�N��c|3��@:�`Q�u���?s#33�4�1K�g�']@g�t�g��&�S`hWm��3�\B����C"�	���81��_�
A�/�4��/�7k �B�W8C?2�� ��� S��4�0�3�� o�=�,�����5ǟ�[����,�I+`������A���>6�jq+ -_������]�s�����������C��U��#Æ��\����O�����M��C(�Cw�j��T�O�D@�+/z�B��( ��7���C�Y������������r�I*�����ڿ	�B���L� �`)��AC�u�g�%�;����v�^C(�B�������"���Ī/J$C�$��ÿ������NA�	�!�7B���?Aw�tJJ3�E����_�T�X����Bv�<�2���"�Dͪ��J��'i�Ϝ����M�A���B�#�C�xA�V��)���C�y��)�����C�8�X`��߄�� [� �������3��� i�^�p��������� ��� /�!S�Hw� ����y������ +=2a�_�q��ÅTD_F�ILTES`i�[3 Է��P��</ /'/9/K/]/o/�/�/ �/6��/�/�/??�,?>?P?b?t?�YSH�IFTMENU [1jWm<�|%� �?�t�?�?O�?�?EO O.O{OROdO�O�O�O��O�O�O�O/__	�LIVE/SNA�P#Svsfli�v�~A_��PI�ON &�U^PdRmenuz___�_�_��r�5G�kΉ��9M�OG�l�~�złZ�Ddm��a<ۀ ��P�$WAIT�DINEND  a�U��#bxfOK-�N�oOUT�o�hS�o�iTIM�e���lGo}�o2{�oz��oz�o�hRELE��.��hTM^{d=�xc_ACTWP-����h_DATA n΅�%�_B��6��rRDIS�P�~��$XVRao�9n�$ZABC_�GRP 1p[k ,2J��=Qa�pVSPT q9m\.�Ԗ
�Z�_���Z)�?�އDCS�CH`r#�����I-Pbs[o!۟����؊MPCF_�G 1t���Q0 O O����u��p�{pK� 	?�t��o`�  ?���2?�k�1�?�ɾ�����4/6��u��D5Oy���C��?�����<� ���>%��6�����u=�!�����ί�>����dن�����˿� � 8��h�Ca��.�~:��1５#����۸���&�  �2�H�Vπ��,�>���0V�h��� �`v�����_CYLINuD�w(� �d� ,(  *E߀V��B��fߣߊ� ��������?� �� D�+�=�z�ߞ���� ����g���@�'�`��v����̞�2x �� �=���?���	��-=��`���zA��SPHE_RE 2y%���� �*����X�k FX��|�� ��///ewT/ �x/_/q/�/��/�/l�/��ZZ�v �f