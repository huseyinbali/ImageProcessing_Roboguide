��   K�A��*SYST�EM*��V9.1�0214 8/�21/2020 A 	  ����CELL_G�RP_T   �� $'FRA�ME $M�OUNT_LOC�CCF_METH�OD  $C�PY_SRC_I�DX_PLATF?RM_OFSCt�DIM_ $BA{SE{ FSETC���AUX_OR�DER   ��XYZ_MAgP �� ��LENGTH�T�TCH_GP_M�~ a AUTORA�IL_��$$�CLASS  O�����D���DVERSIO�N  �VIRTUA�L-9LOOR� G��DD<x$?������kn,  1 <DwX< y�����C�����	/��Z�Zm//�/_/p�/�/�/$ �/��/	?';�$MNU�>A\"�  <��Z9��|���йh0c15���4�
����5!D����࿤oC����0 �?/�?'�?�?�?�? �?!OO)OWO=OOO�O sO�O�O�O�O�O_�O�_A_'_�;5NUM  ����w92�TOOLC?\ �
Y8&,�TP3��E.���P�Q&�TS ;_]_o5_oCo)o[o yo_oqo�o�o�o�o�o �o-%Gu[ }������V�V y�[