��   v��A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@��&�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	�=@&USRVI| 1  < `��R*�R��QPRIƍm� t1�PTR�IP�"m�$$C�LASP ��)�a��R��R `\ �SI�	g�  �aIR�Ts1	o`'2 L1���L1���R	 �,��?����a1`�b�d~a���a��y`� � ����
 ��a�o�o1CU �oz���� �c�
��.�@�R� �v���������Џ� q���*�<�N�`�� ��������̟ޟm�� �&�8�J�\�n����� ����ȯگ�{��"� 4�F�X�j����������Ŀֿ���`/TPTX������/�` sȄ��$/softpa�rt/genli�nk?help=�/md/tpmenu.dg���Ϩ� ���υ�����&�8� J���n߀ߒߤ߶��� W������"�4�F�X� ��|����������+�a�f�f�c �($p�-����T�?�x���a�a��c���c����l���cT��a�dh�h��2�h�	f���������`���`�  ���f ep���h#h�F�d��g�Xc�B 1~)hR \ �_� REG VED]����wholemo�d.htm�	si�ngl	dou�b trip�8brows Q�����u� ��//@/����dev.slh�/3� 1�,	t�/ _�/;/i/??/?�/�S?e?w?�?�?�?� H`�?�? OO$O6O`HOZOlO~O�F @�? �O�O�O�O�O_�F�	 �?�?;_M___q_�_�_ �_�_�_�_�_oo%o 7oIo[omooM'�o�o �o�o�o�o+= Oas����� ����?>�P�b�t� ��������Ώ���O� ����L�^�_'_� ������ş����� 6�1�C�U�~�y����� Ư��ӯ�o���-� ?�Q�c�u��������� Ͽ����)�;�M� _�-��ϬϾ������� ��*�<�7�`�r�A� Sߨߺ�q���i���� �!�J�E�W�i��� �����������"�� /���O�I�w������� ��������+= Oas������ �,>Pbt ���߼���/ /�����^/Y/k/}/ �/�/�/�/�/�/�/? 6?1?C?U?~?y?�?Y� �?�?�?�?�?	OO-O ?OQOcOuO�O�O�O�O �O�O�O__�R_d_ v_�_�_�_�_�_�_�_ �o*o�_o`oro�j��$UI_TOP�MENU 1�K`�aR �
d�a*Q)*default5_�]*leve�l0 * [	 �o�0�o'r�tpio[23]��8tpst[1�[x)w9�o	�=�h58E01_l�.png��6m�enu5�y�p�1!3�z��z	�4���q��]��������� ̏ޏ)Rr���+�=��O�a���prim�=�page,1422,1h����� şן����1�C��U�g���|�class,5p�����ɯhۯ�����13��@*�<�N�`�r���|�53������ҿ���
��|�8��1�C�U� g�y����ϯ���������"Y�`�a�o/��m�!ηq�Y��avtyxl}Tfqmf[0n�l�	��c[164[w��59[x�qG�y�&�tC8�|�29�� o�%�1���{��m�� !�����0�B���f��x���������o���80��'9K~���2P����� \��'9K� �����������1��/$/6/H/Z/�U�|�ainedi'ߑ/�/�/�/�/P��config=single&|�wintp���/$? 6?H?Z?!Z�a�h?�? �e�?���?�?�?O O+O=OOO�?[O�O�O �O�O�O�O�O_a�%_ L_^_p_�_�_�_U��_ �_�_ oo$o�_HoZo lo~o�o�o1o�o�o�o �o 2�oVhz ���?���
� �.��@�d�v����� ����M�����*� <�ˏ`�r���������^��;�M�sc���;���s�� �}����e�u��X��@�F7 L���`��t꒯4�j�X�6e�u7������Ͽ������27��G�Y�k�}Ϗ�� 0�s���������!�1�M�_�q߃� ��T����������� ��7�I�[�m���� ����������!�����6(�]�o��������$��746������)t<ϯ\�5	TPTX[209©|Dw24§J��
�w18��� ����02��A#��[	�tv`�Rx\L�u10�1��5S:�$treeOview3��3��&dual=o'81,26,4� O/a/s/2�/�/�/�/ �/�/�/?'?9?K?]?$o?��;/&�3$/6$ ���?�?�?
?#O5OGO@YOkO}O�?�? "2�?8"2K��O�O_�O���1�?�E��g_y_�_�y6_��edit�� >_P_�_�_o��/�� �_�Cooo�o�oB�o �o��oA�o� +=Oas��o� ������(�9� ��Q�x���������ҏ O����,�>�P�ߏ t���������Ο]��� ��(�:�L�^�ퟂ� ������ʯܯk� �� $�6�H�Z��l����� ��ƿؿ�y�� �2� D�V�h����Ϟϰ��� ���ϕo�o��o@ߧ E�c�u߇ߙ߽߬��� ��O����)�<�M�_� q���W�������� �&�8���\�n����� ����E�������" 4��Xj|��� �S��0B �fx����O ��//,/>/P/� t/�/�/�/�/�/]/�/ ??(?:?L?��߂? 1ߦ?���?�?�?�? O$O5OGO�?SO}O�O �O�O�O�O�O�O��2_ D_V_h_z_�_�_�/�_ �_�_�_
oo�_@oRo dovo�o�o)o�o�o�o �o*�oN`r ���7���� �&��J�\�n����� ����E�ڏ����"� 4�ÏX�j�|������� a?s?蟗?�sO_/� A�S�e�w�������� �������,�=�O� a�#_������ο�� =��(�:�L�^�pς� Ϧϸ������� ߏ� $�6�H�Z�l�~�ߐ� ������������2� D�V�h�z������ ������
����@�R� d�v�����)����������ƚԔ*d?efault%���*level8��ٯw���? �tpst[1]��	�y�tpi�o[23���u����J\me�nu7_l.pn5g_|13���5�{�y4�u6���//'/9/K/ ]/���/�/�/�/�/�/ j/�/?#?5?G?Y?k?~�"prim=|�page,74,1p?�?�?�?�?�?�"��6class,13�?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_B_T_0f_x_{?�218�?�_@�_�_�_�__B6o�9oKo]ooo�o`�$�UI_USERV?IEW 1֑֑�R 
���o��o�o[m�o'9K]  �����l�� �#�5��oB�T�f�� ����ŏ׏鏌��� 1�C�U�g�
������� ��ӟ~�����v�?� Q�c�u���*�����ϯ �󯖯�)�;�M�_�~
�*zoomr�ZOOMIN� q��ؿ���� �ÿ D�V�h�zό�/ϰ����������Z*max�res��MAXRES��	ߧ�p߂ߔ� �߸�[����� ��$� ��H�Z�l�~��;ߡ� ����3���� �2�D� V���z���������e� ����
.��;Q _�������� *<N`� ����w��/ o8/J/\/n/�/#/�/ �/�/�/�/�/?"?4? F?X?/i?w?�?�/�? �?�?�?OO�?BOTO fOxO�O-O�O�O�O�O �O�?__'_�Ob_t_ �_�_�_M_�_�_�_o o(o�_Lo^opo�o�o 7a