��  	c4�A��*SYST�EM*��V9.1�0214 8/�21/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP6fBI�IZ@!�LRM_RECO�"  � ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� ."��!_I�F� � 
$_ENABL@C#T� P dC#U5K�!CMA�B �"�
� �OG�f 0CUR�R_D1P $Q3LI�N@S1I4$C$AU�SOd�APPI�NFOEQ/ 9�L A ?1�5�/ H �7�9EQUIP �2�0NAM� ���2_OVR�?$VERSI� �� PCOUPLE�,   $�!PPV1CES C G�1�!�PR0�2	� � $SOF�T�T_IDBTOTAL_EQ� �Q1]@NO`BU SPI_INDE]�uEXBSCREE�N_�4BSIG��0O%KW@PK�_FI0	$�THKY�GPAN�EhD � DUMMY1d�D�!U�4 Q!RG1R�
� � $TIT1d ��� 7Td7TP� 7TP7T55V65VU75V85V95W05W�>W�A7URWQ7UfW1*pW1zW1�W1�W �6P!SBN_CF��!�0$!J� ; 
2�1_CMN�T�$FLAG�S]�CHE"�$Nb_OPT�2p��(CELLSE�TUP  `f�0HO�0 PRZ1}%{cMACRO�bOREPR�hD0D+`t@��b{�eHM �MN�B
1�UT�OB U��0 9DEVIMC4STI�0�� �P@13��`BQdf"V�AL�#ISP_UsNI�#p_DOv<7IyFR_F�@K%�D13�;A�c�C_�WA?t�a�zOFFu_@N�DEL�x�LF0q�A�qr?1q�p�C?�`�Ab�E�C#�s�ATB�t��d�MO� �sE' � [M�s���2�REV�BI�LF��1XI� %�R�  � OD�}`j�$NO`M�+��b�x�/�"u�� ����!�X�@Dd p =E RD_Eb��?$FSSB�&W`�KBD_SE2uAUG� G�2 "_��B�� V�t:5`ׁ�QC ��a_ED|u � � C2���`S�p�4%$<l �t$OP�@QB9�qy�_OK���0, P_C� y��dh��U �`LACI�!��a���� FqCOM9M� �0$D��ϑ��@�pX��OR BI�GALLOW�� (KD2�2�@V�AR5�d!�AB e`BqL[@S � ,K�JqM�H`S�pZ@M_�O]z���CFnd X�0GR@���M�NFLIx���;@UIRE�x84�"� SWIT=$�/0_No`S�"CFzd0M� �#PEED��!�%`(���p3`J3tV�&$�E�..p`L��ELBOF� �m�� m�p/0��CP�� F�B����1��r@1oJ1E_y_T>!�Բ�`��g���G�� �0WARNMxp�d�%`�V`wNST� COR-�rFLTR�T�RAT T�`� $ACCqM�� R�>r$ORI�.&6ӧRT�SFg WCHGV0I�p�QT��PA�I{�T��!��� � ��#@a���HDR�B��2�BJ; �CѪ�3�4�5�6*�7�8�9>����x@�2 @� TRQ��$%f��ր�׍��_U���ѡ�Oc <� �����Ȩ3�2��LLEC�M�-�MULTI�V4�"$��A
2q�CH�ILD>�
1��z@T}_1b  4� STY2�b4�=@��)24����@��� |9$��T�A�0I`�E��eTO���E��EXT���ᗑ8�B��22�0>�
�@��1b.'��r}!�A�K�  �" K�/%�a��R���?s!>�O�!M��;A�֗�qM�� 	�  =��I�" L�0[��� R�pA��$JO�BB�����`���IGI�# dӀ�����R�-'r��A�ҧ��_�M��b$ tӀF�L6�BNG�A��TBA� ϑ�!��
/1��À�0���R0�P�/p ����%�@|��Bq@W�
2JW�S_RH�CZJZ�T_zJ?�D/5C��	�ӧ��@��Rd&� ����ǯ�r�GӨg@NHANC��$LG/��a2qӐ� ـ@��A�p� ���aR��>$x��?#3DB�?#RA�c?#AZt@�(.�����`gFCT����_F�L�`�SM��!I�+ lA�%` �` ���$ /�/����[�a���M�0\��`��أHK���AEs@͐�!�"WJ��N� S'�I��_'  . II��2�(p�STD_�C�t�1Q��USTJڒU�)#�0U[�m%?IO1��� q_Up�q�* \��=�AORzsBp;�d]��`O6  RSY�G�0�q>EUp��H`G��� {@]�DBPXW�ORK�+��$�SKP_�pAqfa�u�0�TR�p , �=�`����Z �m�OD3��a _C`"�;b�C� �GPL:c�a�tőS�D��G�Bb����P�.�� )DB�!�-,|B APR��
I�Ja3��. /�u���.�� �LUY/b_tS���0�_���P�C�1�_�TENEG�]� 2�_�S6P�RE.��R3H �$C��.$L�c/$USނz )kI3NE�7A_D1%�ROyp�������q0bc7 T@zfPA���?RETURNxb��MMR"U��I�C�RG`EWM�0�SIGNZ�A ��|�e� 0$P'��1$P� m�2��`��`tm�pD�Ip �'�Bd.a	r�GO_AW ���04ؑB1m@CSd�(�KCYI�4���`1w�squ�|t2vz2�vN��}��E]sDEV�IS` 5 P �$��RB��I�wPk��vI_BYȧ��p�TQ�tHN{DG�Q6 H4��1�w��$DSBLC��O��vG@��I�_qL��7/�F@]�fd�FB���FERa@8����t]s���8> �i�T1?���MCS@솀�FD ���[2H� W��EE���%F���λtSLAd��09  ��INP^��]��`�]q��:P +8�S��0x�^���^�,���FI�2���� ���A	AWl���'NTV�㜒V~���7SKI�#TE����0a���T1J_�#;29_�PD�SAF�T��_SV�EXCL�U�῰�D6@L�l �Yք��3�HI�_V
0\2PPLY��@0«�G�����_M�L%��pVRFY�_�C��M��IOC�UC_� ���O�p��LS�`V�&T%4�A1��s���@aPdE&�gp�AU��NFT�u��uZ��pm�ACHD�O���^�6��AFC CPl���TD�4P~�� �� �;�P@T�ѡ0,@_ ���|�N��N=� <Y���T���?� ���{�SGN��=;
$�`�a >aR0I�3�g@ _BM�|_B]�ANNUN�P@~��ÅuC.@�`�/�ɢ�� �����2E�FC@I�R>p�$1F���4OT�`{�@&TD�(RQ<�#QmJ�-Mb�NI�R?��4��6�A��R�DAYCLOAD�tT-��'S5#Q�EFF�_AXI��@�P�QO3O�йS�@_RwTRQ��A D1�t	`��Q,@ ��!EVp�Ӓ���@�0}��0��{��MP�E{� BV������$s��DU�`���.�BCAB��C���P�NS"�+0ID�W�R���V!� V�wVq_���V �DI� ��4D� 1$V�`SEm�TQj�}�'���D�^E_ln�$�VE� � SW���[a���2��A��OH��)�3PP��%�IR�1Bu@p�&���b���� ]�w3W�O � W��vM����C�0��cp��RQ�DWF�MSw0��A�X,���$�LIFE �@����-Q��N�������Co���CB0LqN]a�f��OV0HEQ�NSUP�T���"�@_oS�1_��Gq�Z�
W�
B1�0�#��@�k2XZ_ LQVY2�C9`T_@D``��N�����J�! >�_� ��F� �4�E `�pCACqH,�\�]SIZ(�T ���bN�UFFI� ���@(Td��'S6#Q�1DMp0��F 8��KEYoIMAG�cTM,a�V#��a�^�hB1�OOCVIE�aG�2� L��H���?� �	��D� PH��6�ST'�!C"D��K$PK$-�K$��K EMAILK�u`[��0^��FAUL�RI�28sc�C� COU�0iA��0T`�1J< �$�#�S�m�ITW�BUFp��p(�t�0�0n B�$�t�C�����"�3� SAV-5�"����H7@@��P44�
`�N�a_� 5LЉ9OTgb+���P�P�:���7#AXC����X� T��a3_G��
m@YN�_N� K <\�D��uPb�M�M8�jH TL�F~`$�`��DIزE�@`��aLY���G1��&�G�Da:AF����baM��`A�#�3C_^`�`Knd�@^DQ��R��E�(ADSPl�BPC�KIM:3 �C�A��A��U�Gd meڠ� IP��C7�3�DTH���B�ЙTaa�CHSEC�CB#SC	�"�PV���Z`�P�3�Tp��NVk�AG�S�T�F� F����0d�C5@�1aSC8���u�CMER��Q�FBCMP��~@E�T;� N�FU� DU� ́�`����CD�IYP�0�#m���`NOu�=�O�� �pzbL�xds�P�zbEC"��e
��2�!�uc�0� PH *�aL��_c�q�1f�� ,�'��dD��f"��f-Ѡ�f���f��f7�i8B�i9�j���hz1zU1z1(z15z1BzU1Oz1\z1iz2wz�2{z2z2(z2�5z2Bz2Oz2\z2*iz3wz3z3{zU3(z35z3Bz3Oz�3\z3iz4wr�EXT��=�QB\h@@%@�e@C��e�0�FDR��RT� VW��2�򁑇R��REM��Fq��O�VM�C��A��TR�OV��DT80КMXߜIN��: Ϛ��'IND���
�F@�0@G�1d�ِ9 r��D��ِRIV԰�&��GEAR�AI%O��K��$�N5@���������� %�Z_�MCM� ���Fve UR3bS ,�a�1? 9 P?����?�E@,����1`v�T�j��P�1��RI^e����#ETUP2_� U -��#TDGP0��$Ti��Z�T��qa�"BACBV QTD��"eD)_J%��8�c0@ѰIFI:�0@0`�`�Ь�PT���LUI6$W �� (� URt�1@@�2MA�P� ����I��u$(�Sܰ?x4��Jb@CO|0�3VR�T$���x$SHO8�ѱ��#ASSjP�18(IPQ�BG_�����s��s��(s��5sF�ORC�"7��DAkTA��X�"FUס�1:B��2:ALOG����Y |*�N;AV�0�(�X�����S�"&$VgISI[�.BSC�4�SE�t�7�VB�O
r���Bò�A�Z֯$PO,�IE���FMR2s�Z ��i`f⁑ s@�օ�������ǖ� ��堒_wqX���I#T_ֱSd��ME�j��|�DGCLF;�D7GDYd�LD�H�!5
?�ѡMcp8#�[��� T�sFS�07$\ P2����sC�0$EX_������1�0�PE��53�5��G�Q��g] ��0bSW5}O��DEBUG��L]�GRc��U�S�BKU`O1�p  PO�Ј�t��"`G�t�Ms�LOO,�3��SM�E<2|���& _E ^ y��TERM��9_��� ORISA��y`��cp�SM_`@�]���a������ b���~�UP"c�3 -�D�^(����f _>�Gk
}�EL�TO�!>B�PFIGf?AנS�`b�`$UFRfB�${`�� Ne�OT���PTAiP���N;STT@PAT^Qi��PTHJ&aL`Ep9 d2U`�ARTU0��� U1�">AREL<Ac1SHFTPR?A3__�R/`Ic% ) $8�b.႐8S�S�2SHId+��U�b O1AYLO .P�1 A��j����e[PERV p�� �$��T@A��Ȱ+%̫�ȰRC��eAScYM3A�e?AWJ�$� �E$�/[)�OaU$T@ A3��&IaPS��Q�ORT@�M��/����d���t��� �16�H9Os���e �˶,s�i`OC���$OP^��A�cFv���a�i@��2R0R�S"OU�Se�R�5m8K���e$PWR]�IM�5"R_H3(*И ?AUD$�kS�Voc1SDfH�$�HdE!@ADDR
C�H��G7A,A%Ap"�p@F��ag H2�S�PFѝ�dE��dEs�dE(sSE��H��`H�SY`MN�h�W�@0��"QebaOL�/SW�{0R�\f��AC�RO����ND_�C/Szb��4�QROUP�S2_��
Ғ�11�q��:S�DY3  DY��EXpDY(pDY��⊒AC���SAVE�D?W�SOUG�C��gi $��@0_D)�x��j«BPRM_
�}~�HTTP_z`�H�aj (;`OB�JB�%B��$C�L�E�0a�`k �� 4��6�_�TĽ�XbS0�3��KR�L�9HITCOU����G�LS�j0Xbb�`$�f�j0ʷk0SS����dJQUERY_�FLA�C_ _WE�BSOCI��HW�cq�+�l_@� IONCPU�R*�Ov ma��K�0pzD/q�D/q~ǂ�IOLN���m 82�R��i��$SL��$INoPUT_��$�0�~xPy� mZpS)L�P+�nep{�u`�tB#�uB"NAIO�P�F_AS��o��Q$��B��qN�Yр�2��ksM�ts�H�YB�5���A�pUOP��p `�pS�C�@��%���,�}��0P�3��0s���,������I�P_ME\��q �X�pIP,@�Rւ_!NP��`*�G2B��O��BSP���P��F�BG�Q�-�M<!��r l �TA4�3`As�TI���%�� ��_�OPS^�BU��ID�Ўbs����x0��;a-���� sD�r?�r�S��pNҘ���ӕ�IRCA_�CN� t ��Ji�pCY�@EA ��C��q��31�#���@z"���!DAY_<����NTVA�����u��r#��u�SCA��u�CLO᎑j����@��u��ڔ$��N_R0Cβ򐎒c�6�v�r��^3%����'b�����Pi��� �2u �����wp��\�'b\�LAB��z��Ѐ�UNIбn�	 ITYl�.�0E"��R; G���x�r��R_URLЀ$A�AEN|�k�*��0��CT�AT_U#� ��Jp��yр$�_%E�pRk�.���AS��q8�J�aC�F�L��K��P
W�r�
��UJR�%z ��J`F��(����D�£$J7S%�J�8��7&�h�����7����8�ɭ�APHMI�Q����D���J7J8"�L_�KE��  ��KQpLMܑ { <٠XR�p$p��WATCH_VA��A�ű#fFIEL��"Cy��2Ҳ�| �
��V�G-1��CTpܰ������LGɳ�}� !�LG_SIZRdv��հ�����p��FD��I ���ة����������� d3��V��V��pV��@V���V�K!G�� _� _CM�������AF�!�����А4(������������p��� �I��
���0��������RSU��  (.p�L�N���"~_��`DE��E�r!�s���S��0L���DAU��EA�PQp44����GH52X��pBOO~YA� C��ʀIT�c��� �R9E4�SCR��|c��D�PKr,QMARGI�q�;�v�S4He�d�qS8c�rWC��q���JGM�MgNCH���qFN(�b�K����	UF�ܯ�FWD�HL.STP�
V���X����RS?H� ��C�~"�� w�U�Q�v�Ȩ���G�	PPO �"2�� ��	�EX�TUI�I ;���;�8bZ#�Z#� ���R��P# r#N�A�3ANA�rA1��AI���D�� �DCSf�lC�#zC�"O�(O�'SK�2�(9S�(ZIGN�Ў�`����4��$DEA|LL"�
��q����i��м�T��$�׀��r
���n2�A����۠lp*s�AV��S1�52�53�1p.�"� �Ђ �Jk�0�$�u�t���Q`�e���:FSTe��R��Y�B\A �$EkFCkK���P�zF�F��#�у L p#�n�8����Co`���d�P�Dtm�}#_ � �Pt��Px��$ S�MCt��� �J`CLD�Pe� �TRQLI0��"�PY>TFL%�iR��QrS��D��rWpLqDrU\TrUORG(��v�R��RESERAV2t�T>s�TIr /S~v�� � 	[UvMTrUSVd�PP^��	�Q+d3fRCLMCAd�_�_SiTp3a�|�MDBG�qͰ��?�$DEBUG�MAS&�_�P���U�uT� |�E�����MFRQV�߈ � ��HR/S_RU�q�A'�yA5��FREQ�����$� ��OVEARt���F��P�7EFI��%�A(��a���c�T� \8�q��$U@%�g?`��PS�0
C�	sC��BcN��s�ScUݐ�a?( �	{�MISCuŊ� d}�ARQA�	f�TBN �� �m!�AX �-��.�EXCES벽��r)M��̱����r �쾱�rSC@ � H"�	�_S��8�P��,�>�.PKɴ��rد�N �eB_��FL�IC�DB QUI[RE�MO��O��pv�QL�@Mȵ� �P��E����AbF�aND��q�ހ�{��r��؄�D���IN�AUT4��RSM����+0N$bn�j��PSTḺ� 4n٠LOCFRI��vEEX�ANG�"ܲq�aODA�e�b�p|����MF�� �Cv7I�BA �Eq�o�ΨfSUP�EwqFX�;�IGG � �`�Cn�(�C� �Da�br\B��^@ɨ^@�ئ���P��7�qTI�vл��Po�M+��b�� t9�MD6���) D�� O�XaL�H����O�DIA��P�>�W�iO��1�O�D��)p/�t�)`ހ� m�CU��V��#`�qՁ�O\_�`y�� �`��CC��`rr��B �P �J���P���KE�^���-$B8+p��@ND2ZbZ��P�2_TX�DXT�RA�#|�lb�E�L�O��ހ�k����	 ��u�ǲ�ƪ�%��RR2�u�� �.����A0a d�$CALI�o�Gt�!��2�0RIN�����<$R��SW0�_d,�lcABCJ�D�_Jb����pC�_Ju3W�
Q�1SP��$���pPQ�x�3w�̱�@�p��Jlc���R�(aOu1IMl`�rCSKP_Z�Ի��#��	J���rQ��������_AZ/b��I��ELZ1��ZaOCMaP��q�q��RT�a�t��1��В��1ї��{ ��Z��SM�GY'�zdJGPS�CLN�
�SPH_@0�p7��㓰�p��ORTER+���� R��_� Q6@A\ �SC�r'�DI_���2[3U��DF{�H�LWN�VELPQIqN�Bf q�_BL� �ry��ѳqJi�~�����MECH�2lbwq#IN
�q���ǲ���]�q ��@_�p �����/��`��1���?�ՀDHN�~�:����0$V������{!$��'qrA�+$O1.PR������H �$BE�LZ��g�_ACC�E� �la� I�RC_(��a�PNyT�q;C$PSN�
CRL{���XS�� �?�� �G��	�"3�ؠQ�_�1l�IO"u�p�_MG�sDDl(�rFW�3P(�����}D}E�PPABN�RO��EE_�1��PP��1�a���{��$USE_���#P.+pCTR�$Y�~ Z.a �AYN�pAm 6&��f�6!M�aұ�"�fOk�
c$INC �������'���ENC�L��r�X��� INCBI���%)���NTi��N�T23_L�r�#L!O]�r09pI\�� 6R���p���0����yC���&MOSIq���߰O!s�rPER�CH  ��7q�  y7��3�2zd�o� g� %&N��A��5L$�ӻ����%��:�F36TRK��AAY���3��HA�WELC��z暁�"�`MOM }"����P̰����acC���DU���DS_BCKLSH_C��E�`X68p�>#�s�C�"ZM!�CLALM�$�a�@ �5UCHK���Z�GLRTY��A��$��Q'�_f�M4_UM�c�VC�cz��Sp7LMTt�_Lj b��Tv��WE�]�P�[�P ��U��нc�2 d�8PC�1�8H��&�p��UCMC��z~C�N_	�N��f��S	F��9V "��'�pTa��eXhCAT�^SHf�	�~�&yQ�A��&����ɗ�mPAL�T�"_P�UrC_�Ѐ��OFm0��_CqtbUJaGJ�d�esW�OGrg>�TORQU �� K3hI��c2��r_W�EHD��m�t^��ud�uI�{I
�IdF0��q��I���v�VC� 0����j�1�p�n��0�v�JRK�p�������DB��Mt����M��_DL^�2GRV�t�^�dՁH_��Ӄ"��COS/�|�/�LN ��R�s�Y�^ T���T� &���~�D�ЅZM�c6ՁMY[�Θ;�I�C���THET0#5N�K23d�X\�C�B�CBXC��AS�C�&�Q�^Q���SB^o�)�GTS���C{�Kq��:s��<����$DU_P�7�ʢ��٧��Q�1_�4cqNE��K oT��-�< �A�:�pC�!�,�,�LPH/���%�Ss���~���������������:�V�\�VQ�N t�V��V���V��V��V��V
ȻVֹH\�u�{�s���a�Ȑ�H��H��H���HȻHֹOM�OR\�O�r�O��O��UO��O��O��OȻO��F�>���~����O�SPBALANgCE_ޑ��LE��H_�SP��o����~��ҍ�PFULC�����⍕��1����UTO_ZPbUTg1T2^�2NAQ �� ~���A������AT	@OA��p�INSEG�<1R�EV��<0�!DIF�2E	1���?�1��%@OB��%Q���G2��p� LQ݄LCHW3AR�%"ABAq�E���<0ސU!���SX�UAPdt�3�?S��� 
u��q��%RO�Bm0CR�2��ib � �C�_]rT� � x $�WEIGHR p�$M���tpIR!0I9F
!�LAGC""bqSC"��C"BIL)cOD�@?0ST� "P��%P  | �`������
� �D!�]q  2�J4D�EBULX�ɠMMY9���N8+s�p$D�1�$� op � �  �DO_� A�� <��rh��$D!0�BB: N�#�_!0D _O2P ��� %�PT�� �!�QT��� TgICK-�T1� %j�@sNm0M�	m0R�@D!=�=��� PROMPR#E~/� $IR�p�B!hP��0"MAI�ڀ}!T"�_# ����^AV R�CO�DwFUJ ID�_�0'%�����G_�SUFF&� h9!��DO�0���< �GR#=� e$�q$=�|%=�%�q�e$�� ���H�_�FIv9�#OR�DB ��36�b�"B!� $ZD�T.%�0_��4{ *��L_NA�s52�DEF_I E852�Q4�I�S`�}3��5�IS�@�`���3�O4D�a�4�abSDQ�(�B�4wD�pO�� LOCKE+q_#�`���1e"_ UMd% 52e$}3e$�5e$�2q" gCp%`3q$�4q"Q�F �1|#H�^q|%52|%}3 |#�GUa(8P�4H�1�� WFHEU<C� 1TE0Q��� LOMB�__RzW0VIS�=�ITYAoqO>CA_FRIN�SF�SI�1�Q�RpH�W{�W3�W�X!W�[倩V��_i�!EAS�"�q�Tp�@��V4�Y5�Y6�ORMULA_�I+q�G%7� �h �7�COEFF_OW��d$W��GqS ��CA���_GR�� � � �$<@��
XGTM�/G't<E]DCA|E�R��T%D$4� � M G�LL�$@S/�g_SV�4�x$hV� ����d� � �rSETU�3MEA�D b� _�"�� � �p�� � �` �� �A�":2sA0AD�bA�Q�";��@�1�@G����RE�C�!�2SK_���s� P��1_USERz�j���p,𾔙�z�VEL>� ��,�����=�I0��w�MT8CFG����  u��Oc�NORE�� ���-��� 4 ��s^�d�XYZ��#�������_ERR�� ��ep6� �c\�}��Ҁ�� BUFINDX�1���PRt� H��CU\�d���1Ӄ���!$���10����W��Gr� � $SI�`�P ��Ɲ�VO
����OB�JE��ADJU���AY9p���DJ�OU� 5���C!.�"=��T��y�8��x��DIR}���p�������DYNb$����TR�5�R�QH�B 4��OPWOR�� �,� S�YSBU*�2�SO!P���q�U���1P<@߂4�PA���X6�_�2�OPz U4��(��t�e�IM�AGo���q�SIM��IN`\���?RGOVRD��%���g�Pi��������@( C׵d�L:@BY���> �PMC_E0���N*�M±�1��2��SL����{ ���OVSL��S:RDEX�1�0K�2c���a_��cǬ  ��cì mÂ�}Ȫ�ÁC��70���Ƿ�_ZER �*��s��G� @"���~�O/ RI���
����ɠ�����'�L����T`�W ATUS�p�C_T����O�B+pY�B���3�.�0��� D�e�N� LҾ��M��!��o��XES���һ҆���1�����R�UP:��0��1PX�y�b��3�ǂ���PG텳>��$SUBA�~���AA��JMPWA�IT��r�Y�LOWp/�^�' CVF��vc�\�R���q�C�C��R��i��IG�NR_PL�DB�TBW P�1d�BW� ���U*��IG�L��Ic�TNLND����R֡5B�PN��E�PEED��T�HADOWW b����ES�M�b�+�P0SP]D��� L��Ar�0Q0m�/�{�UN �dy���R�м�LY0���K�'�PH_P�K����RETRcIE��i�y!0����FI�� �x:����� 2����DBGLV��LO�GSIZ��1KT�y�U�s2D8� �_[TX�EM�`Cn����X ARR.R+�C�HECK��1��)P��p�c������LE�4pPA#@T���C�O��P��p��bAR%"���#�1�'�O� 0��`ATT ���x�%X ��1Ɵ�UX���PL�,  $��/QS�WITCHT��aW��AS���SL�LBp�� �$BAv�D
C2�BCAM�������#J5L���6�|_KNOW�����U=�AD��`x�D���)PAYLOA��@%#_��.'�.'�Z+#L�AA�q�0L�CL_ʐ !@�pg"�Ӂt$˲�&F�)Cgpb*�e$�`�Ib(Ripb'{�~$Bd7`ʑJ���!_Jl!:��֑ANDz�U�`
4l"�!(�"aPL�?AL_ �`x�Pѐ����PC>�D*#�E=��J3036�{ T�`PDCK��22�CO�p_AL3PHC3�3BEБsa�C?U<��b��� �� �.�$/D_�1+*2U$D�pAR���H�5FC�TI�A41I51I6>�MOM��=C]CJC]CWC�Bp�AD=C�FJC\�FWCPUB�RbD �EJC�EWB�@30ʑ�q�  � MO"L� �T����� e$PI ����3��0'&Y��J)*&YI2[I@[INS�D S�V�V�ޠ2p������1�HIGo 1�q�j��Vj�q������V�S�X���Y��q�SAMP�Я�:d�W;c8q�3 �pia ʐS�Œxd��fj��0 �i@Œߠ�:@�e/02��H��cIN�l/0 c�h�k�dq��jx�d�{2{GAMM�eS|U�A�$GET�Rd��3�D�4҂
$60�IBR���IL�$HI:�_����Œ�v�Eѐ�xA�~�p�vLW�}�v�|�y��v�2�V�51C��CHKhİ��q�x>I_` �ޔ.2�8.1�e|�uC�ޔ�F{�33 ��$e8 1��I��RCH_D��Ɩ�RNs�8���LE@���R����8Ѐ��MSWFL���AS;CR�100{�. xd39]��gʐ=@�ixq�j���PI3AVMETHO�æ���V��AX$���X4�p�ERI��:d3�fsR�� 5	�Q�0FHWt;ac��c��(�L�;a=�OOP�a֑S��a֑APP��F� W�x�c�&�cRT��2�O0j��0�������DR 1��%��D��ѪNPѢRA֟ MG�OSV�	Q�P; CUR�C��GRO7���S�_SA�ܴ5���NO�0C�����45��t �?6/H/TX����zP�X�UϸCDOi�A�r dyes��e�X��W� �X3�/��k#���D��T� � ��YQL$S�!�g��S�"6A9��K���!������!_�C���M_Wd���C�����?�M���ˇ ��21~�AL�T�K�� PM&�R� �}�R��YWE�S$��L3 X!EШ4Cү4CҶ4C�W4���pN��sf��J/0X��O�3.1Z�ո P{�T� ���M��z�w���������@4@����� �C�1_Z� |v1��5�]I�� JC��WC5�6J���PJ�uu 9 p������Y s�P��P�MON_QU?` �� 8� QCO�U��QTH_�H�O~�:�HYSES�:�UE%�+�� ]OX�  ��P#���uV�RUN_TOʱ���O�R
P� �P! ��C����I�NDE�ROGR�A��J��2C�NEg_NO���IT�A���g�INFO���C b��������OI��� (SLEQ�V"�U" ���A�OSU��� =4� ENABqҁ�PTION
�ERVE�R~�Q�VwGCF_� @.�J �.1����pR³��T_EwDIT��� �R�R��K�A�S�qE�psNUAUTQ�	COPY�A�P*�Q]�M�qN48M��PRUTR ;N� OUC�Q$G�����RGADJn��� hv0X_��AI���п�пW��P����S��rN^0_CYCq��/RGNS[�s�=��LGOZ��PNYQ__FREQ�BW�`��VP!SIZn[�L�AœG!�XC�`�UCcRE�p��[�IF@Q���NACa%�$_}GœSTATUv�<œy�MAILAb�1x�!
�5�LAST�!��1"$ELEM_�� �\�iFEASIl3�nbg�Z�2�� >�96���`�pI�����G"�Q=� ��n2AB$U�0E���PV�!�6�BAS�2�5�r�AU8�P�PJ�$�1�7RM�@Rh3Ł���3`���P�r�!�4 ��$"S�~�	E2 2� �c���d +F�2*G�2"Э`���28VGW�DOU�����r�"$P �@�)G�RID��U�BAR�S�WTYm "OT�O����� t�_"�$!��B�DO��\�� � ����P�OR���C���CSReV� )TVDIS�T_�P4PFT�PPW�P�PW4NY5NY6NY7�NY82Q�Fbr_�~r�$VALU�3�(�+4��Q\��C !h^����C�!%���AN'��R�!���T")1TOTAL_X�$l06bPW=#I�A>KdREGENIj^b��X�8��=�� f �cTR�3�"Ia_S+��g^`��V���b��2E�# �?�(2�� ncV_H�@DA ��`pS_YY���a&�S8�AR �2� }�IG_SE6�ȷ`R�%_���dC_��F$CMm�f�wrD�Eh�?p�rI]�Z�vsPsq!�F��HA{NC&�� pA�j�"d#qINT�1P��F}���MAsSK퓸0OVR���� �<�!Ł�Gy��	��Q�E�d�OJ6�k>�F�PSLGHp�Q� \ 1�b%Z��$�3`� S���$�qUY�y����c��ZQ�Us�TE��@�' (�aJV�Q��q#IL_Mp$�Vt2����TQ ���R�0C���VB�CP��P_�J�Z�Mq�V�1p�V1~�2��2�~�3��3~�4��4 ~�� ��<�����;IN�VIB0�J��7��>�2:�2F�3*:�3F�4:�4F��� Y�r�U��gP
�tP���'��PL� TOR$��IN��u��5����T $�MC_FC�X�B�LC�B��u)`M��1I�s*�rC ��)���r��KEEP_H/NADD#�!e��0o�C�ѳ����A$�����O�d�>"��`����w��REM��@���!�Bµٱ޸U�$�e��HPWD  ;e�SBM�q�@?COLLAB"��Ph��'a�" IT' ��INO)�FCAqLh�
���� ,���FLnб1$SY�N���M��Ccr�~�`UP_DLY��=�r�DELA���!Z�"Y �AD �.��QSKIPG�� 	�
P��O��˂K���P_����Ƕ��� ��#ٖ#�gP"�tP "ځP"ڎP"ڛP"ڨPz"�9��J2R *���dX�0TJ#�� ��)1�Ѭa�����a���RDCaw�� %�� R��R�!�8=��-DRGE� W3�{BFLG�0��sSW{	-DSPC���!UM_����2T�H2NuA��� 1�  ���|�A[ � D��x�x]�02_PC����S���1Q L10�_Co"����q ���JPٰ7��6K�@+��� �.�NE����N���b\r�3����p����DE�SIG��JEVL1b��1��k��10ٰ_DS�K�j��`C;11��� lV���0����iI�AT��� �AS'J N$	C��
���HOME�4 ���2��� ���� 2D����3���gy����� ��4�����,>�5���as����S ���6����@�//&/8/V7���[/m//�/�/�/J'8����/�/�/? ?�2? ��S)�������1��s`Y�V۰=E�D� T���4L,f�3IO��
II�0:XrOe�_OPE.Cx&b�3�POWE��� �0����8�P/�'c �}�eB�$DSB��GNA�r�%c��C���Q�Sw232�5� ���Z5��׀ICEU�S/cSPE���QP�ARITq$aOPyBQ��RFLOWAp�TR�01b�UJsCqU�@6��QUXT�q|�Q�pERFAC�D�ʰU `J"SC�H�Q� tV��_��@kpc�$�`�`O	M*p��A>�#�p%��UPD<����aPT��0|uEXЙX|S!%�FA?��r��q�a � ���`;b- K�AL$� ��U���]B�a  2�� �S���0�	O� �${�����WGRO�`*dT��(p6fDSPBfJO�G�`�C����AZ�N�������"VK�P_�MIR^a~d�MT3��cAP%����`}t��Sp�`R��
��eBRKHUQ�V��wAXI�1  �b�c�r-b�q9�7e�`B�SOC6f۰N2uD�UMMY16O�7$SV��DE3A�C)F�wK�0�D�pc�OR{ws0N�p|vF�p�w[`OV^eSFN�zRUN�s�rF�v�Q�cUFRA�zTOTLCH�����#OVlt[�[`WP�7� [c���r?p��_�p�� @h�TINV�EG@n1OFS\�C�P�WD�q��q>qXf2�eXpTRr��1�a�E_FD�aM�B_CW���B��B��*��ałˁ?�epV@9Q��P&��írGƇ�hAM�c��VP�F�!�_M݀R_�CS��T$����Q�3T$�HBK�Q�fm�IO�5|�&A��PPA p���������,�&BS�?DVC_DBъ0 ސ�Q�Bސ7�Q������F���3��L�E����+P�`lqU�3P`FCAB�Ё2~㷀8û`� ���O�UX�fSUBCP�[�-�� /��P/Ѯ�ރ��bB��$HW_C@��	P/ы��?�q0�#��P�$UP�t|	��ATTRIh���h`CYC��g�C�AB��cFLTR_2_FI�3�IH��F���PtkCHK�_�SCT�cF_�F1_����FS�A��CHA�}�ֱ�RղRSD���Aq�S�A&@_T�}�.�L��PEM�0��MsTò/��Pò��K��DIAG�URAI�LAC듑�M`L�O"p��Hv_�$P�SNb�2 ��L��P�RߐS}�I���Ctёf�	E�FUN��*QRIN1�}�|00^���Q�S_;`��X����0f���P�f�GCBL���.�A'�#�*�#�DAp��h�.�'�LDyP`p����dCa�����TI�������P$CE_gRIAa�BAF���P�A��~���T2b}�C�S�؁OI����DF_L�0�r�Q��PLM�F^�HRgDYO�af�RG���H���a|0p�/�MULSE�����Qp�$JxzJ�r�w�{FAN_ALMp���WRN��HAR�D�0�VZ0P]R�2����A��e_��fA�U�RȴRTO_SBR&E�O`#���ӓ��;�MPINF�Q��N��Y�RE�G�6NV�Pf3�fD�A@N��FL����$M�Ѕ�`S����P�����CMѐNF�-��1���h��A�v�0$�1$Y �oQb�Q�0�7� ��cEG�0+c�`p+AR=`CHu2�5Rr:T��eAXE�EgROBBjRED&BfWR,� q_�$sCSY�`ep�S��WRI,�>�ST�r@CcPp�pE�D�0G6Rr��;`B� �R��7��2�OTOri��0��ARYBc`4~�2��"t`FI�`~�c$LINK��GTHS�PT_��R�F8Rr|X�YZ�R�9�OFIFZ�S{o8	B@`���/��@�P�FI1�����CXt��Zd_J�A�R�r``����30Rr �@�*!m�b"CFA�e�DUn�Hu3����TUR��X�ӛ%BI�1X� `�J'FL|��a�8 � ��	3ʡ^g� 1��0Kg`M�d�&Qs�����°�pSORQ&�Oa�P(���`O� �1ɐj4��8Ma��~4OVE�1MIPk1��5�5��6_Q�7c��7��4ANڡV�1���1�` �0�k1�5�1�7(E�(E�3OaERla�	B��E,��P��fDAA�P���!�@o�l�o�AX/��Ro�2�� U�EQ��I{��I���J N �J�J$�J��J��J1[ �F/��I/� �I/��I/��I/�Y/� Y/�(Y/�8Y/�HYeQ�YYDEBUڣ$�����I�	ao�wAB�o�m��q3Vb�٢ 
$b�LeʡXg QqXg��XgNXgXg $Xg�Xg���g ��\U�LAB�J5֠�GRO[�J"��K�B_/�MF��s � �v5qK51u�=vAND0��[DL��^A�zw K���� �x01ѝxN�NT��#��pVEL5��4�qm���x9��NA���V�$��ASS ? ����* �*  �_�SI�@��#�ㅆ)�IY�n��(�A�AVM��K 2 �T� 0  �5�䋏������ ���	݀΍�* U��ߏ��!�͌@�L��܁R�������e�BSܿ1  16�� <u���� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲������߸�߱��pMAX/� ����ʓ  d��IN�*��PR_E_EXE;�g��J�!43��T�e�IOgCNV�"<� �&��P��a ;�Ɨ��IO�_�� 1r�P $b�����V���U�?�����$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ�����LARMRECOV ~�!�J����LMDG ����� �LM_IF ��+��ߥ� ��ɯۯ骓���0��B�S�, 
  S�|��������ƿؿ�$�����1��U��g�yϋϝ��NGT�OL  ~� 	? A   ������PPINFO Z� Y��*�8<�N�!�  f�P� ~�?�mߧߑ��ߵ��߀���%��5�[��� �χ������������)�;�M�_�m�P�PLICATIO�N ?����H�Ha�ndlingTo�ol �� 
V�9.10P/30���j�
8834�0����F0����1�028���������7DF1��j���N�onej�FR=Aj� 6w�_ACTIVE�s  ����  ��UTOMOD� �^��ÊCHGAP�ONL� �O�UPLED 1��� 
 2��CUREQ 1]	��  T<<<	����@��<�����Hk�?HTTHKY�A� o���////�/ S/e/w/�/�/�/�/�/ �/�/??+?�?O?a? s?�?�?�?�?�?�?�? OO'O�OKO]OoO�O �O�O�O�O�O�O�O_ #_}_G_Y_k_�_�_�_ �_�_�_�_�_ooyo CoUogo�o�o�o�o�o �o�o�o	u?Q c������� ���q�;�M�_�}� ��������ˏݏ�� �m�7�I�[�y���� ����ǟٟ����i� 3�E�W�u�{������� ïկ����e�/�A�`S�q�w��NTO�����DO_CLE�AN���NM ; �� <_��qσϕϧ�BDSP�DRYRϊHI� ;�@L��%�7�I� [�m�ߑߣߵ������߇MAX~�������	�X��>�PLUGG� ��\�PRC��B9�E=����c�Oh�����SEGF� K ������9�K��%�7�pI�[�����LAP�� ������������	 -?Qcu��TOTAL+�T��_USENU���� ޸��NRGD�ISPMMC��20�C���@@����O������_S�TRING 1
~�
�M� �S�

^_ITwEM1h  n� �������/ /&/8/J/\/n/�/�/�/�/�/�/I/�O SIGNAL�bTryou�t Modei�Inp0Simu�latedmO�ut,<OVE�RR�� = 10�0lIn cy�cl 5mPro?g Abor63m�4Status�k	Heartb�eatgMH �Faul�7�3Aler�9�/�?�?�?O�#O5OGOYOkO}O ��d��v�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ oo�OWOR��dJa �O$oro�o�o�o�o�o �o�o&8J\�n�����~POb�1�pbk��#� 5�G�Y�k�}������� ŏ׏�����1�C�8U�g��rDEV�~�� ����˟ݟ��� %�7�I�[�m���������ǯٯ����PALT�M6�bo�^� p���������ʿܿ�  ��$�6�H�Z�l�~�8�Ϣ�$�GRI�d ��N�����&�8�J� \�n߀ߒߤ߶����� �����"�4�F���� R�M~���X����� ���� ��$�6�H�Z� l�~�������������l�PREG:�# �� ��J\n���� ����"4F�Xj|��-�$A�RG_J`D ?	�������  	]$�&	[�]����')�SBN_?CONFIG� ��$1#2=!!CI�I_SAVE  ��$F!9#�TCE�LLSETUP ��%  OM�E_IO�-�,%MOV_H� �/�/�REP���/�UT_OBACKv!��@"FRA:\� �/F '�`�0C8� �T;?  2�3/07/18 �17:50:04(�?�?�?�?4<��O6OHOZOlO~O�O�$O�O�O�O �O__�O<_N_`_r_ �_�_�_3_�_�_�_o o&o�_Jo\ono�o�o��o�o���  /1_�3_\ATBCK?CTL.TM���o�+=;INI�9�v56%J!0MESSAGV dqF!�>o{ODE_D� Y&�6%�xO���3PwAUS� !��� , 	�� ���,		 �8�"�\�F�X���|� �����֏�����F��t�pTSK  ��}C?I0UPD�T�pbwd���vXWZD_ENBbt2*��STAau�����XIS$ UNT� 2�C!E �� 	 )��� ��4_�D `� ����
���+����:6D�:�s�F��Е��/6�5\�5 [^. 8��a�¯����\����MET��2i��b# P�BZ�A���A���d73�
A�߳A��٭>a�:>ٻ�>p��35ؔ>B��>H�0�S�CRDCFG 1��%1 �^%C"篻�Ϳ߿���<?
QZ)��e� wωϛϭϿ�&���J� ��+�=�O�a�����1GR��������`NA� �	�4��_ED`p1���� 
 �%=-�`EDT-���*��B��b?$� -(3�
"O�&�
��  ����2��#� �G��_���@G����6����3� �+]���̔\��Z�l�����4K��� ����t�&8�\��5�d���@@���(��6� S0/w��/w/��f/���7�//�/C/ ���/C?�/�/2?�/��!8{?���?�f&��?@OV?h?�?�?��9GO�?�O�?i&�pO�O"O04O�OXO��CR���/ __q_ =:_�_�O�O�_�"_����NO_DE�L�ߞ�GE_UN�USE�ߜ�IGALLOW 1���   (*SYSTEM*֣�	$SERV_�GR�k_`�pREG�he$�c֬_`NU�M�j�c�mPMU|`֥LAY��֬PMPAyLap�eCYC1p�Ăc }�`�n%sUL�SU�o�mr�qjc�L;ttBOXOR=I�eCUR_ap�m�PMCNV�f�ap10~�pT4�DLIǐZ|i	*�PROGRAgd?PG_MI�n�F)�AL�u6� �)��BT�_n$FLU?I_RESUw���o��ÄMRvn�`�\�_Β��+�=�O� a�s���������͟ߟ ���'�9�K�]�o� ��������ɯۯ�����#��RLAL_OUT Nk���WD_ABORp�/o��ITR_RT/N  �D��ل�?NONSTO�Я�� 8hCE_RIgA_I,`��������FCFG ����ĨN�_L�IMvb2�� �  � 	��DgϳB<�҄��e�@� VϷ����ϨHa
��ߒ�2�PAn��GP 1��ޥ�n߀ߒ�Q�CO>  C.���f��Qz���߶Ї�Б��U��Р�Ъ�д���������������C����ǀ CѶ���J��G?��HE�PONFIπ��d�G_P�p1;� �U;ծ������������,�d�KPA�US~q1;��� �r.�t�;�b����� ����������0 @fL����6��M��NFO 1v?�� �T���B�̵���5Au�9�	�]�Ǝ�@���K D5�Oy���C����($6��T5+��P�� 8�h�C�a��.~:��1５�ⰍO�ϨG��COLLECT_�a?�x�ǯEN�pp������NDE��?�;c�R1�234567890'�Bya�//&��	HC��C)j/�/y\i/ {/�/z[�/�/?�/�/ ?`?+?=?O?�?s?�? �?�?�?�?�?8OOO 'O�OKO]OoO�O�O�O��O_�O�9��� ��IO !)������_�_ض_�_`WTR6�2"D](�{Y
�O�^o��#o] jt�i_MkOR9�$;� ��HB�!;`�e  �i�o�o�o�o�o�kbbT1�:�%pm,t�?]�]���>q�KFt�
`�R�&�utqtr�C4  A���Ț�x�A����BʤpCd B��d C7  @�r��q�:d�QbZqI#'d}?�s9�(pm����}dZqT_DEFB� {%oR��thPNUSE��s���g��KEY_TBL � ������	
��� !"#�$%&'()*+�,-./(':;<=>?@ABC)��GHIJKLMN�OPQRSTUV�WXYZ[\]^�_`abcdef�ghijklmn�opqrstuv�wxyz{|}~���������������������������������������������������������������������������,��������������������������������������������������������������4Q��L�CKp�ٹ��p�ST�A���t_AUTO�_DOζkv�I�ND�ٞ�R_T1���T23�ݵʳ���TRL(�LE�TE��z�_SCREEN ;ڿkcsc�U�ʰMMENU 1)l� <7�@�� ����F��#�I��� Y�k��������ſ׿ ��6���l�C�UϢ� yϋϱ������� ��� 	�V�-�?�eߞ�u߇� �߽߫�
������R� )�;��_�q���� �������<��%�r� I�[������������� ��&��5nEW �{�����" �X/A�ew�����/)\ʠ_?MANUALo�*��DB'a.b����DB�G_ERRL.�9*֫�Q /�/��/�.L!NUMLKIM���lu
L!�PXWORK 1+֫�/#?5?G?Y?|k?mDBTB_��G ,{-�s�Qst�3QDB_AWA�YT#�QGCP �lr=���"�2_A!L� ٟ�2P"Yn���tlpE(_n  1-�[,p
?POJf@O}O6�6_M�IS֐�;�@�p�CONTIM6���lt��FI�
� CMOTNE�NDt�DRECO�RD 13֫ y��OxsG�O�KQ 9_x{�2w_�_�_�_DX �_�_K_ oo_$o6oHo �_�_~o�_�oo�o�o �o�o�o �oD�oh z���1�U 
��.�@��d���� �����Џ�Q��u� ���N�`�r���󏨟 ���;����&��� J�5�C������ȯ 7��ׯm�"���F�X� j��y����Ŀ3�� ��ϣ���Bϱ�f�տ �ϜϮ���[���S�߀w�,�>�P�b��Ͽ2TOLERENC�4sB�B�0L��L �CSS_CNST_CY 249�Y 	e�B��������� �#�5�G�]�k�}�� ����������������DEVICE ;25�� �6o� ���������������&�O��HNDG�D 6�۬0Cz�9
Q��LS 27Y�8������:��PARAM 8,I�2�5&��ySLAVE �9YE_CFG� :F&d�MC:\��L%0?4d.CSV%@�c�B�A �C	H kkO&/B/
X�&2"_!o/])<\!1@JPя#N.�A�1n_CRC_OUT ;Y���1*_NOCOD�z<,G�SGN� ="UR#M��18-JU�L-23 23:�46�0A:917:�51�~� V�hr9n1&o061��M��Þ�ǧj��1�>�VE�RSION �):V4.2.�11�KEFLOG�IC 1>�� 	�(1@I�!M��2PROG_ENqB Xa=CULS�G� `�2_ACC�LIM�F����|CWRSTJ�NT�G
S���1MO�FLX!2�DINIT� ?��"U�� �FOPTu ?	��F�B
 	Rg575&'P74,Y56-X7-W50QX�4�WR2-T�({_�7
TTO  ]�?�_�6]V�@DEX�Gd�B�� �SPATH ;A):A\�_5o�Go|�HCP_CL?NTID ?�6� �+Ӈo���IAG_GRP {2D� �� 	 D� � D�� D � B��Т��f�f�j�`���o�l�a����%��B��N�C�-BzBp��e`��imp2m7� 7890123�456xq�G�`� � Ao�
A�j{Ad�]���AW�AP���AJ=qAC3w3A<�4z�jL�p�!@��]pA�q���A�����B�4�lf�dX�!
��ru�ppQ�Aj��HAeG�A_��pY��AS�pM�2�F�RA@(� �J���t�J��I��@�p��������@��HL�^�p���������33<���=q@~�R@x�Q�@q�@k��@dz�@]��Vff؏����� ���s>�l��@�e@^J�W
�=@Pv�G�@u@v�7ڐ.{d��v���������S>�M����AR�<(�@�5Ґ/\)@(��@!R�֏ �� $�6��ĭ���ܯ"� 4����V�|�Z����� <�N�������0�B� ̿R��B�`�r5���M�xّe��m>��R���?�33?9���{���m7'Ŭ���6��4�F���L�m@ž�����ڐ␀N�Њ=@V�pAh�����c�= c<��]�>*�H>V�>�3�>���~�m<���<b��a�i�L. �?�� �C�  <(��UX" 4� >��ё��ٝiA吳 ?�el���t����,� �H��8�b���r��z�x����x�?�7���>�(�>!�����=����m��G��G��m�����I��m����i�@��Ҁ�@Q�?L ��Ly�o�g�v\����]p'�@����8����	�gC� �̇�Cu��Zl �<� ���`��&%�18� �����4J�6�<�D5�OL��rC��� >T&U�Q���$�z�	��($6�T��Á�i���x�������=ʝm;��t���9/�aCT_CON?FIG E?i3�eg�%�aSTBF_TTS�G�
UI�#�0�C�A�&�� MAU�@JOJ"M_SW_CFX F�k�  �p�:OCVI�EW� G�-�a���o=?O?a?s?�?�? �B+?�?�?�?�?OO �?>OPObOtO�O�O'O �O�O�O�O__(_�O L_^_p_�_�_�_5_�_ �_�_ oo$o�_HoZo lo~o�o�o�oCo�o�o �o 2�oVhz0���@,RC�#{��"!L�~���A��0�e�T����$SBL�_FAULT �I�z 8��GPMS�K�'��L TDIAOG J\)�!���1�UD1�: 6789012345�p"1�j'�uP&/O�a�s����� ����͟ߟ���'� 9�K�]�o�����y���
>���F&TREC	P���
���%��� =�:�L�^�p������� ��ʿܿ� ��$�6πH�Zρ�������7U�MP_OPTIO1N� ����TR�"�#:����PME�%���Y_TEMP  È�3BȞ �1��A.��UNI�� �%1��&YN_B�RK K?6EDITOR����
���_ԠENT 1�L�y  ,&�MAI��TLO�G T1��e�&GPAR���߫����2��0�&OMAY�[���F��߇� ��� u���J�����
IRVWAI�����&-BCKE�DT- ��/����PICKSIM_���[���y���o"� x������������� 3WiP�t�������~�MGDI_STAD�� !1�y�NC71M�+ �`�r��
��d�����/ !/3/E/W/i/{/�/�/ �/�/�/�/�/??/? A?S?��j?|?�?�?�9 ��?�?�?�?
OO.O @OROdOvO�O�O�O�O �O�O�O__*_<_�: c?m__�_�_�?�_�_ �_�_o!o3oEoWoio {o�o�o�o�o�o�o�o /A[_ew� ��_������ +�=�O�a�s������� ��͏ߏ���'�9� SA�o��������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�K�]�g�y� ��A�����ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� C�U�_�q߃ߕ߯��� ��������%�7�I� [�m��������� �����!�3�M�W�i� {����߱��������� /ASew� ������ +E�Oas���� ����//'/9/ K/]/o/�/�/�/�/�/ �/�/�/?#?=/?Y? k?}?���?�?�?�? �?OO1OCOUOgOyO �O�O�O�O�O�O�O	_ _5?G?Q_c_u_�_�? �_�_�_�_�_oo)o ;oMo_oqo�o�o�o�o �o�o�o�_?_I [m�_���� ���!�3�E�W�i� {�������ÏՏ��� ��7A�S�e�w�� ������џ����� +�=�O�a�s������� ��ͯ߯���/�� K�]�o��������ɿ ۿ����#�5�G�Y� k�}Ϗϡϳ������� ���'�9�C�U�g�� ���߯���������	� �-�?�Q�c�u��� �����������1� ;�M�_�q��ߕ����� ������%7I [m����� ��)�3EWi ��������� ////A/S/e/w/�/ �/�/�/�/�/�/?! +?=?O?a?{m?�?�? �?�?�?�?OO'O9O KO]OoO�O�O�O�O�O �O�O�O?_5_G_Y_ s?�?�_�_�_�_�_�_ �_oo1oCoUogoyo �o�o�o�o�o�o�o_ #_-?Qc}_�� �������)� ;�M�_�q��������� ˏݏ�i%�7�I� [�u�������ǟٟ ����!�3�E�W�i� {�������ïկ��� ��/�A�S�m�w��� ������ѿ����� +�=�O�a�sυϗϩ� �����������'�9� K�e�[߁ߓߥ߷��� �������#�5�G�Y� k�}���������� ���1�C���o�y� ��������������	 -?Qcu�� �������) ;Mg�q���� ���//%/7/I/ [/m//�/�/�/�/�/ �/?!?3?E?_i? {?�?�?�?�?�?�?�? OO/OAOSOeOwO�O �O�O�O�O�O�/__ +_=_W?I_s_�_�_�_ �_�_�_�_oo'o9o Ko]ooo�o�o�o�o�o �o�O�o#5O_a_ k}������ ���1�C�U�g�y� ��������ӏ�o�o	� �-�?�Yc�u����� ����ϟ����)� ;�M�_�q��������� ˯E�����%�7�Q� [�m��������ǿٿ ����!�3�E�W�i� {ύϟϱ�������� ��/�I�S�e�w߉� �߭߿��������� +�=�O�a�s���� ����������'�A� 7�]�o����������� ������#5GY�k}������ ��$ENETMO�DE 1NB��  �������� R�ROR_PROG %�
%��an�<TABLE  �L������<SEV_NUM� 
  �� <_AUT�O_ENB  �(9_NO! �O� " W *�Y �Y �Y 	�Y  +X r/�/�/�2$FLTR/0&H�IS���++_A�LM 1P� e���Y,��+�/�2?D?V?h?z?�?�/_\�8   �W!��:� TCP_V_ER !�
!Y��?$EXTLOGo_REQ�&�))�#CSIZ,ODST�KIIG%� BT�OL  ��Dz��"�A D_BWD�0�@�&�A#�C�DI�A QB���C��KST�EP�O�O� �@OP�_DOkO�FAC�TORY_TUN��'d3YDR_GR�P 1R�	�!d �	�?�_{P�*�u���RH�B ��2 ���� �e9 �����V{S�_�]{PB����B�A�C���B���Aן�BM��@�[A��K�A�B���&A���A?I��B� �[ �_WoBo{ofo�o�o�o��o  @�:A|=@9q��o���
 F�5Wx&b�`��A����o�	2�o�o\G��]��  �qA��`�3�3�r�33�]@UUT�z@�`�pj$�>u.�>*���<����]E�� F@ �p&���]J��NJk��I'PKHu���IP�sF!�=��]?�  j���9�<9��896C'�6<,5����~���=�����a�� ��_&���#tF�EATURE �SB��@"�Handling�Tool 	����English� Diction�ary�4D S�t��ard	��A�nalog I/�O@�I�gle S�hift\�uto� Softwar�e Update���matic B�ackup���g�round Ed�it��Came�raW�F[�Cnr�RndIm���o�mmon cal�ib UI��n�͑�Monito�r&�tr�Rel�iabp��DHC�P�]�ata A�cquis5�^�iagnos��T�x��ocument �VieweA�`�u�al Check Safety!�~�hanced!�4���sʠFrސ��xt. DIO �1�fi��&�end.��Err@�L��B�J�sA�rR�1� �@��FCTN Me�nu�v\���TPw In��fac���GigE��εƐ�p Mask Ekxc��g#�HT���Proxy Sv�ˤ�igh-Spe��Ski�Ŧ�~5�mmunic��7ons<�ur�����s�X���conne�ct 2s�ncr��stru#�qʚ��e��۠J���KA�REL Cmd.� L �ua���R�un-Ti"�Enyv�Ȅ�el +���s��S/W�LicenseݣʬX��Book(Sys�tem)�MAC�ROs,3�/Of'fsew�V�H5����q�[�MR:�6���MechStop�t����V�iS�s���ax��T�����odq�witch�ߚӡ�y.{��Optm,��filʬ��g�i�V�ulti-T���Г�PCM fun�Ǣ�o��ޢ��^��RegiK�rW���riàF����U�Num Sel��|� � AdjuG���=�s�N�tatu���f�Ū�RDM �Robot �scgove)���ea���"�Freq An;lyW�Rem��5��n7�����Serv�o5���SNPX� b�x�SN��C�li¡%t�Libr(�E�� ��W �o0�t��ssag����0 ��n���0�/I���MILI�B��P Fir�m���P��Acc<ǐϛTPTXm��elnn����j�޲orquq�imGula?��bu��PaѱƐZ�(�&��ev.���ri�۠:USB poort �iPL��aà�R EVN�T��nexcept����������VC�rR�I���V@��o"�%Wz+S8 sSC4�/SGE�/��%UI�Web Pl}� >i�'4������x�ZDT ApplP��&?|7�Grid��pla�yv=� ���7Rf".�7��6���/Y�-10�iA/8L�?A�larm Cau�se/��ed*�A�scii�<�Losadʠ:JUplP@2�l�7�Gu=�rO2�BP��Ֆycp���0��蠕�RA� ��9�NRTJ�O}n�e Hel���漿������1tr�;�ROS Ethj
�t�BeW7iR�$�2D Pk;�uVI�m+�Fd�� �^ns�p���Q�64MB� DRAM�O�SFsRO�_ېellW�F�shao gcK�de��p�2ltyp�As'�ԗ�B��D�.�maiܠ;�JT�qV�R7��FL!PSup�c��� pL���cro~���W�4x��&��auestz&�rtڡ���/�3D�L}|�Q���Ty,K���l Bui��n��/APLC��uV�Z��/CGl��CR�G#��$D��@�R�L�S[��%BUw��%K�і��!TA���Bp�,يE�TCB���ʏ��/��^�T�C��v��%��TCEHǟٖ"�ؗV�����/��F�H�����G:���n�������H¯��IA߯�ޯ��LN���M��D���HD�����N���P��H������RR���Sڿ�����W.�@Ǣ��$gVGFf�x�P2Z� ��2��ǂϔ�B�ϔ�	D�ϔ�Fr�����"7TUT��01J�\�y2f�\�TBGG��ކ�rain��UI�*ЦUHMI��r pConU2�8���af{ ��R�v�VKAREL���_TP� �e� �R9�0�B�o�f�x�� ������������5� ,�>�k�b�t������� ��������1(: g^p����� �� -$6cZ l������� �)/ /2/_/V/h/�/ �/�/�/�/�/�/�/%? ?.?[?R?d?�?�?�? �?�?�?�?�?!OO*O WONO`O�O�O�O�O�O �O�O�O__&_S_J_ \_�_�_�_�_�_�_�_ �_oo"oOoFoXo�o |o�o�o�o�o�o�o KBT�x� �������� G�>�P�}�t������� ׏Ώ�����C�:� L�y�p�������ӟʟ ܟ	� ��?�6�H�u� l�~�����ϯƯد� ���;�2�D�q�h�z� ����˿¿Կ���
� 7�.�@�m�d�vψϚ� �Ͼ��������3�*� <�i�`�r߄ߖ��ߺ� �������/�&�8�e� \�n��������� ����+�"�4�a�X�j� |��������������� '0]Tfx� ������# ,YPbt��� ����//(/U/ L/^/p/�/�/�/�/�/ �/�/??$?Q?H?Z? l?~?�?�?�?�?�?�? OO OMODOVOhOzO �O�O�O�O�O�O_
_ _I_@_R_d_v_�_�_ �_�_�_�_oooEo <oNo`oro�o�o�o�o �o�oA8J \n������ ���=�4�F�X�j� ������͏ď֏��� �9�0�B�T�f����� ��ɟ��ҟ�����5� ,�>�P�b�������ů ��ί����1�(�:� L�^�����������ʿ ��� �-�$�6�H�Z� ��~ϐϽϴ������� ��)� �2�D�V߃�z� �߹߰���������%� �.�@�R��v��� ���������!��*� <�N�{�r��������� ������&8J wn�������  H5�52��21R�7850J6{14ATUP)�545)6VC�AMCRIdU�IF)28eNR�E52XR63�SCHDOC�V�CSU86�9)04EIOC��4R69XEgSETAWJ7W�R68MASK^PRXY}7OCO(3A! �(3`&J6'53��H�(LCHH&O�PLGA0x&MH�CRI&S�'MCS�@0$'554MD�SW!7k'OPk'M�PRl&��(0(PCM|R0g7! 4l� �'51L51�8�0LPRS'69�`&FRDdFRE�QMCN93�(SNBA��'SHLBFM'G�8�2(HTC@TMsIL�TPA�oTPTXYFEL�6�� �8J9�5�TUTl'95�`&UEV&UEC�H&UFRdVCC� XO�&VIPdFC;SC�FCSG���IWEB@HT�T@R6��HCG�_WIGGWIPGS��VRCdFDGk'H�7�R66LR7�'R�8R53�76U8�82x&R�*4�W�664R64NVD&R6�'9 �XX�9 �D0+gF~h�CLIP8KCMS���`@STY$WT�O@NN`&ORS��&M�8OL�hEN�DLWS�hFV�R�V3D$X{P�BV�FAPL�A�PVl&CCG@C�CR�&CDWCD�L�VCSB�CS�K,6CT{GCTB�HV�p�hC(F�p�xC�<WTC|�ppwTCv�wTC&CTE��9�|wTE�9�0WTUF�xF�hG�xGx�
$�H$�IF��$��GWCTM�hM�M�xUN$�P��P�xR�x��hTS�xW8��VV�GFP�P2 WP2��6e�\�B\�D\�F6|VP��VT���VTB�wV�I�HWGV�P՗K$WV _V��)�;�M�_�q� ��������˯ݯ�� �%�7�I�[�m���� ����ǿٿ����!� 3�E�W�i�{ύϟϱ� ����������/�A� S�e�w߉ߛ߭߿��� ������+�=�O�a� s����������� ��'�9�K�]�o��� �������������� #5GYk}�� �����1 CUgy���� ���	//-/?/Q/ c/u/�/�/�/�/�/�/ �/??)?;?M?_?q? �?�?�?�?�?�?�?O O%O7OIO[OmOO�O �O�O�O�O�O�O_!_ 3_E_W_i_{_�_�_�_ �_�_�_�_oo/oAo Soeowo�o�o�o�o�o �o�o+=Oa s������� ��'�9�K�]�o����������ɏۏ�  H55Ȕp�����R78�{50	�J614	��ATU�?�545z9�6	�VCAM	�wCRI��UIF9��28��NRE�5�2x�R63�SC�H	�DOCV��C�SU�8699�0^H�EIOCɛ4(��R69x�ESET�Y�w�J7w�R68��MASK	�PR�XY��7	�OCOBy�3Y�(���8�3ت[J67�53(�H��LCH��OPLGzY�0��MHCR��]Sw�MCSX�0��{55H�MDSWٻv�OP�MPR�t�(�08�PCM���R07˅�H���(�5�1h�51x�0h�P�RSx�69تFR�D��FREQ�M�CN	�938�SN�BAٛ�SHLB�	�M7��ȼ28�H{TCX�TMIL��(�TPAH�TPT�Xy�EL�ʅ�(�8�'�%��J95��T�UT�95تUE�Vx�UEC��UF]R��VCCX�O��wVIP��CSC�ڧCSGȚ�I	�W�EBX�HTTX�R�6ל��CG��IG޷�IPGS	�RC���DG�H7'�R[66h�R7g�Rv̷R53h�68h�2j��R6�4��66H�wR64�NVDx�R6����h��������D0��FVCLI�g�CMSH�� X��STY��TOX�N]NتORS��M�̻OL�END�L�g�S�FVRH�Vs3D�짛PBV��wAPLH�APV�wCCGX�CCRx��CDg�CDL(�C�SB�CSK�CT��CTB�� ��C8�5 ,C��TCب�5 �TC�TC�x�CTE��� �T�E�� ��TF,FJ�G,G�-�,H�,�I�E0�,��CTM��Mx,M�N�,P�H<P,R,�TSr,W�=(�VGFKP2X�P2��5@(L�B(LD(LF��VP�W;VT��@(�VT�B�V�IHw�V5��KK��V���_ 1_C_U_g_y_�_�_�_ �_�_�_�_	oo-o?o Qocouo�o�o�o�o�o �o�o);M_ q������� ��%�7�I�[�m�� ������Ǐُ���� !�3�E�W�i�{����� ��ß՟�����/� A�S�e�w��������� ѯ�����+�=�O� a�s���������Ϳ߿ ���'�9�K�]�o� �ϓϥϷ��������� �#�5�G�Y�k�}ߏ� �߳����������� 1�C�U�g�y���� ��������	��-�?� Q�c�u����������� ����);M_ q������� %7I[m �������/ !/3/E/W/i/{/�/�/ �/�/�/�/�/??/? A?S?e?w?�?�?�?�? �?�?�?OO+O=OOO aOsO�O�O�O�O�O�O �O__'_9_K_]_o_ �_�_�_�_�_�_�_�_ o#o5oGoYoko}o�o �o�o�o�o�o�o 1CUgy��� ����	��-�?� Q�c�u���������Ϗ���STD~�LANG� � �2�D�V�h�z��� ����ԟ���
�� .�@�R�d�v������� ��Я�����*�<� N�`�r���������̿ ޿���&�8�J�\� nπϒϤ϶������� ���"�4�F�X�j�|߸�ߠ߲�RBT�OPTN����������#�5�G�Y�k�DPN ������������ ��%�7�I�[�m�� �������������� !3EWi{�� �����/ ASew���� ���*�/1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? OO)O;OMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/AS ew������ ���+�=�O�a�s� ��������͏ߏ�� �'�9�K�]�o����� ����ɟ۟����#� 5�G�Y�k�}������� ůׯ�����1�C� U�g�y���������ӿ ���	��-�?�Q�c� uχϙϫϽ������� ��)�;�M�_�q߃� �ߧ߹��������� %�7�I�[�m���� �����������!�3� E�W�i�{��������� ������/ASe�h�������99��$F�EAT_ADD �?	���~  	� %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�? �?OO+O=OOOaOsO �O�O�O�O�O�O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_�_o#o 5oGoYoko}o�o�o�o �o�o�o�o1C Ugy����� ��	��-�?�Q�c� u���������Ϗ�� ��)�;�M�_�q��� ������˟ݟ��� %�7�I�[�m������ ��ǯٯ����!�3� E�W�i�{�������ÿ տ�����/�A�S� e�wωϛϭϿ���������DEMO �S   �N�D�V߃�zߌ� �߰����������� I�@�R��v���� ����������E�<� N�{�r����������� ����
A8Jw n������� =4Fsj| ������// 9/0/B/o/f/x/�/�/ �/�/�/�/�/?5?,? >?k?b?t?�?�?�?�? �?�?�?O1O(O:OgO ^OpO�O�O�O�O�O�O �O _-_$_6_c_Z_l_ �_�_�_�_�_�_�_�_ )o o2o_oVoho�o�o �o�o�o�o�o�o% .[Rd���� ����!��*�W� N�`�������Ï��̏ �����&�S�J�\� ����������ȟ�� ��"�O�F�X���|� ������įޯ��� �K�B�T���x����� ����ڿ����G� >�P�}�tφϳϪϼ� �������C�:�L� y�p߂߯ߦ߸����� 	� ��?�6�H�u�l� ~����������� �;�2�D�q�h�z��� ����������
7 .@mdv��� ����3*< i`r����� ��///&/8/e/\/ n/�/�/�/�/�/�/�/ �/+?"?4?a?X?j?�? �?�?�?�?�?�?�?'O O0O]OTOfO�O�O�O �O�O�O�O�O#__,_ Y_P_b_�_�_�_�_�_ �_�_�_oo(oUoLo ^o�o�o�o�o�o�o�o �o$QHZ� ~������� � �M�D�V���z��� ����ݏԏ��
�� I�@�R��v������� ٟП����E�<� N�{�r�������կ̯ ޯ���A�8�J�w� n�������ѿȿڿ� ���=�4�F�s�j�|� �Ϡ����������� 9�0�B�o�f�xߒߜ� �����������5�,� >�k�b�t������ �������1�(�:�g� ^�p������������� �� -$6cZl �������� ) 2_Vh�� ������%// ./[/R/d/~/�/�/�/ �/�/�/�/!??*?W? N?`?z?�?�?�?�?�? �?�?OO&OSOJO\O vO�O�O�O�O�O�O�O __"_O_F_X_r_|_ �_�_�_�_�_�_oo oKoBoTonoxo�o�o �o�o�o�oG >Pjt���� �����C�:�L� f�p�������ӏʏ܏ 	� ��?�6�H�b�l� ������ϟƟ؟��� �;�2�D�^�h����� ��˯¯ԯ���
�7� .�@�Z�d�������ǿ ��п�����3�*�<� V�`ύτϖ��Ϻ��� �����/�&�8�R�\� �߀ߒ߿߶������� ��+�"�4�N�X��|� ������������'� �0�J�T���x����� ����������#, FP}t���� ���(BL yp������ �//$/>/H/u/l/ ~/�/�/�/�/�/�/? ? ?:?D?q?h?z?�? �?�?�?�?�?O
OO 6O@OmOdOvO�O�O�O��O�O�O__2]  )XH_Z_l_~_ �_�_�_�_�_�_�_o  o2oDoVohozo�o�o �o�o�o�o�o
. @Rdv���� �����*�<�N� `�r���������̏ޏ ����&�8�J�\�n� ��������ȟڟ��� �"�4�F�X�j�|��� ����į֯����� 0�B�T�f�x������� ��ҿ�����,�>� P�b�tφϘϪϼ��� ������(�:�L�^� p߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�h�z����� ����������
. @Rdv���� ���*<N `r������ �//&/8/J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П�����*�<�N� `�r���������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ�����������>0�  1�6� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~������ �� �2�D�V�h�z� ������ԏ���
� �.�@�R�d�v����� ����П�����*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������(�:� L�^�p����������� ���� $6HZ l~������ � 2DVhz �������
/ /./@/R/d/v/�/�/ �/�/�/�/�/??*? <?N?`?r?�?�?�?�? �?�?�?OO&O8OJO \OnO�O�O�O�O�O�O �O�O_"_4_F_X_j_ |_�_�_�_�_�_�_�_ oo0oBoTofoxo�o �o�o�o�o�o�o ,>Pbt��� ������(�:� L�^�p���������ʏ ܏� ��$�6�H�Z� l�~�������Ɵ؟� ��� �2�D�V�h�z� ������¯ԯ���
� �.�@�R�d�v����� ����п�����*� <�N�`�rτϖϨϺπ��������&�5�:�-�P�b�t߆ߘ� �߼���������(� :�L�^�p����� ������ ��$�6�H� Z�l�~����������� ���� 2DVh z������� 
.@Rdv� ������// */</N/`/r/�/�/�/ �/�/�/�/??&?8? J?\?n?�?�?�?�?�? �?�?�?O"O4OFOXO jO|O�O�O�O�O�O�O �O__0_B_T_f_x_ �_�_�_�_�_�_�_o o,o>oPoboto�o�o �o�o�o�o�o( :L^p���� ��� ��$�6�H� Z�l�~�������Ə؏ ���� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X� j�|ߎߠ߲������� ����0�B�T�f�x� ������������� �,�>�P�b�t����� ����������( :L^p���� ��� $6H Zl~����� ��/ /2/D/V/h/ z/�/�/�/�/�/�/�/ 
??.?@?R?d?v?�? �?�?�?�?�?�?OO *O<ONO`OrO�O�O�O �O�O�O�O__&_8Y��$FEAT_D�EMOIN  V=T�hP�=PPT_INDEX][lQ��PPILECOM�P T�����QkRKU�PS�ETUP2 U��U�R�  �N �Q�S_AP2�BCK 1V�Y  �)9Xok%�_:o=P�P(oeo ;U�_�o o�oDo�o�o zo�o3E�oi�o ��.�R��� ��A��N�w���� *���я`������+� ��O�ޏs������8� ͟\�ڟ���'���K� ]�쟁������F�ۯ j������5�įY�� f������B�׿�x� Ϝ�1�C�ҿg����� ��,���P���t���� ��?���c�u�ߙ�(� ����^��߂��)�� M���q� �~��6��� Z������%���I�[� ��������D���h�@����
3�Y�PP�_� 2�P*.V1R:���*��`�����n PC�|��FR6:�"4�X�T|P| �y�_PI����*.Fq/��	��<,�`/�STMk/�/"�/�-O/�/�H�/?�'�?�/�/i?�GIF s?�?�%�?F?X?�?�JPG�?!O�%O�?�?qO�
JS{O�O���7C�OOO%
Ja�vaScript�O�?CS�O(_�&_��O %Casc�ading St�yle Shee�tsT_��
ARGNAME.DT�_
��� \�_U_�A�T��_�_�PDISP	*�_���To�_�Q�Na\oo
TPEI?NS.XML�o�_�:\�o]o�QCus�tom Tool�bar�oiPAS�SWORDSo��FRS:\#�oD`�Password Configd ���<���� +�=��a������&� ��J�ߏn������9� ȏ2�o�����"���ɟ X��|��#���G�֟ k������0�ůT��� �������C�U��y� �����>�ӿb����� ��-ϼ�Q��Jχ�� ��:�����p�ߔ�)� ;���_��σ��$߹� H���l�����7��� [�m��ߑ� ����V� ��z�����E���i� ��b���.���R����� ����AS��w �*<�`��� +�O�s�� 8��n/�'/� �]/��//z/�/F/ �/j/�/?�/5?�/Y? k?�/�??�?B?T?�? x?O�?OCO�?gO�? �O�O,O�OPO�O�O�O _�O?_�O�Ou__�_ (_�_�_^_�_�_o)o �_Mo�_qo�oo�o6o �oZolo�o%�o [�o��D� h���3��W�� ������@����v� ���/�A�Џe�􏉟 ��*���N��r��������$FILE_�DGBCK 1V������� < �)�
SUMMARY�.DG#�ϜMD�:W���ېDi�ag Summa�ry����
CONSLOG��p���ۯ����Conso?le log���	TPACCN��v�%^�����TP� Account�in=���FR6�:IPKDMP.'ZIPϿӘ
� ������Except�ion$�ջ��ME?MCHECK����􆯧�/�Memory Data�Ͼ�� l�)��RIPE��ϒ�'߶��%�� Pac�ket L<���L��$�e���STA�T!��߯� �%C�Statuys��`�	FTP�������1�mment TBD4��`� >I)ETHERNEy��f��w�瑱Ethe�rnL�3�figu�raCϫ��DCSVRF(�� �9������ verif�y all<���M�.c��DIFF�1��)���=�S�di�ff��t�f���CHG01������C��X��kv�- 	29� 2���hz3p���K ��rVTRND?IAG.LSw(�:���� Op�e��N� ��nos�tic���)�VDEV�DA�T������V�is�Devic9e�+IMG���./@/�/<�k$Imsagw/+UP �ES/�/FRS�:\?\=��Up�dates Li�st\?��� FL?EXEVEN��/��/�?���1 UI�F EvO�O���,��t)
PSRBWLD.CMO�ϜG2#O^?0�PS�_ROBOWEL<U���:GIG�ϾO��?�O��GigE��(O��N�A�)}�AHADOW�O��O�Oi_��Sha�dow Chan�ge�����a�~)RRCMERRa_�F_X_�_���PCFG Errorq �tail�_ MA��m�CMSGLIB�_�_�_so�B6e���|0ico+a�)_`ZD�O�o\o��o��ZDPad�o l )RNOT�I��o�ow��N?otific�� F�AG���՟� ���(���L��p��� ���5�ʏ܏k� ��� $�6�ŏZ��~���� ��C�؟g������2� ��V�h��������¯ Q��u�
����@�ϯ d�󯈿��)���M�� ����ϧ�<�N�ݿr� ϖ�%ϣ���[���� �&ߵ�J���n߀�� ��3�����i��ߍ�"� ��/�X���|���� A���e������0��� T�f�������=��� ��s���,>��b ����'�K�� ��:�Gp� �#��Y�}/ $/�H/�l/~//�/ 1/�/U/�/�/�/ ?�/ D?V?�/z?	?�?�??? �?c?�?
O�?.O�?RO �?_O�OO�O;O�O�O qO_�O*_<_�O`_�O �_�_%_�_I_�_m_�_ o�_8o�_\ono�_�o !o�o�oWo�o{o" �oF�oj�ow�/ �S�����B� T��x������=�ҏ�a������,���$�FILE_FRS�PRT  ��������A�MDONLY� 1VU�� �
 �)MD:�_VDAEXTP.ZZZ3�䏻�ʛ�6%NO �Back fil�e ���S�6) �����@�	�M�v��� ��)���Я_������ *���N�ݯr������ 7�̿[�ٿϑ�&ϵ� J�\�뿀�Ϥ϶�E� ��i���ߟ�4���X� ��eߎ�߲�A����� w���0�B���f�������E�VISBC�Ks�]���*.V�D����U�FR:�\��ION\DA�TA\��w�U��Vision VD��!�[�m���� {��D�����z��� 3E��i���. �R����A �Rw�*�� `��/��O/� s/�/@/�/8/�/\/�/ ?�/'?�/K?]?�/�?�?�?4?F?�?;�LU�I_CONFIG7 WU����;� $ �3x�{ U�=OOOaOsO�O�O�I%@|x�?�O�O�O_ _'\�OJ_\_n_�_�_ )_�_�_�_�_�_o�_ 4oFoXojo|o�o%o�o �o�o�o�o�o0B Tfx�!��� ����,�>�P�b� t��������Ώ��� ���(�:�L�^�p��� �����ʟܟ��� $�6�H�Z�l������ ��Ưدꯁ�� �2� D�V�h���������¿ Կ�}�
��.�@�R� d����ϚϬϾ����� y���*�<�N�`��� �ߖߨߺ�����u�� �&�8�J���[��� �����_������"� 4�F���j�|������� ��[�����0B ��fx����W ��,>�b t����S�� //(/:/�^/p/�/ �/�/=/�/�/�/ ?? $?�/H?Z?l?~?�?�? 9?�?�?�?�?O O�? DOVOhOzO�O�O5O�O �O�O�O
__�O@_R_ d_v_�_�_1_�_�_�_ �_oo�_<oNo`oro(�o�o&h�`x�o�c��$FLUI_D�ATA X�����a�)a�dRESULT� 2Y�ep ��T�/wi�zard/gui�ded/step�s/Expert �o?Qcu���������S�kip Gpan�ce and F�inish Setup�D�V�h�z� ������ԏ���&hW �`.)`�e>!�0 �2`!���c�aA��ps �������ԟ��� 
��.�@�R��2oy� ��������ӯ���	� �-�?�Q�)e�)cA��3�E�W�g�rip *pu�ۿ����#�5� G�Y�k�}Ϗϡ�`��� ��������1�C�U� g�yߋߝ�\�n�����䤿b�g�%pTimeUS/DST�� ?�Q�c�u������������
�Enable��(�:�L�^� p���������������
 �b�a���������#�24*�� �����1 C��y���� ���	//-/?/Q/�"4F\�$qRegionT/�/�/ ??+?=?O?a?s?�?��?�AmericaϿ�?�?�?OO +O=OOOaOsO�O�O�)aym//�O�/�/#sditor�O7_I_ [_m__�_�_�_�_�_��_� Touch Panel  S� (recommenp)�_>oPobo to�o�o�o�o�o�o�o�L��O�O5�O	_Racces�?�� �������,��>���Conne�ct to NetworkM����� ����̏ޏ����&�(8�J��H�^ 9+�=S!_PInt?roduct�/� ����*�<�N�`�r� �����Ϻ�̯ޯ�� �&�8�J�\�n������� ��w�����Y>VSafet�A$� 6�H�Z�l�~ϐϢϴ� �����ϩ�� �2�D� V�h�zߌߞ߰����� ���߷�ɿ��[� k�}���������� ����1�C��g�y� ��������������	-?[(�5��-�Q���� �"4FXj| �M������/ /0/B/T/f/x/�/�/ [m�/�??,? >?P?b?t?�?�?�?�? �?�?��?O(O:OLO ^OpO�O�O�O�O�O�O �O�/_�/3_�/Z_l_ ~_�_�_�_�_�_�_�_ o o2oDoU_hozo�o �o�o�o�o�o�o
 .@�Oa#_�G_� ������*�<� N�`�r�����Uo��̏ ޏ����&�8�J�\� n�����Q��uן� ���"�4�F�X�j�|� ������į֯诧�� �0�B�T�f�x����� ����ҿ俣��ǟ)� ;���b�tφϘϪϼ� ��������(�:��� ^�p߂ߔߦ߸����� �� ��$�6���?�� c��Oϴ��������� � �2�D�V�h�z��� K߰���������
 .@Rdv�G�� k����*< N`r����� ���//&/8/J/\/ n/�/�/�/�/�/�/� ���1?�X?j?|? �?�?�?�?�?�?�?O O0O�TOfOxO�O�O �O�O�O�O�O__,_ >_�/?!?�_E?�_�_ �_�_�_oo(o:oLo ^opo�oAO�o�o�o�o �o $6HZl ~�O_a_s_��_� � �2�D�V�h�z��� ����ԏ�o�
�� .�@�R�d�v������� ��П⟡��'�� N�`�r���������̯ ޯ���&�8�I�\� n���������ȿڿ� ���"�4��U��y� ;��ϲ���������� �0�B�T�f�xߊ�I� ������������,� >�P�b�t��Eϧ�i� ��Ϗ���(�:�L� ^�p������������� �� $6HZl ~�������� ��/��Vhz� ������
// ./��R/d/v/�/�/�/ �/�/�/�/??*?� 3W?�?C�?�?�? �?�?OO&O8OJO\O nO�O?/�O�O�O�O�O �O_"_4_F_X_j_|_ ;?�?_?�_�_�?�_o o0oBoTofoxo�o�o �o�o�o�O�o, >Pbt���� ��_�_�_�_%��_L� ^�p���������ʏ܏ � ��$��oH�Z�l� ~�������Ɵ؟��� � �2����w�9� ����¯ԯ���
�� .�@�R�d�v�5����� ��п�����*�<� N�`�rτ�C�U�g��� ������&�8�J�\� n߀ߒߤ߶��߇��� ���"�4�F�X�j�|� ������������ ���B�T�f�x����� ����������, =�Pbt���� ���(��I �m/������ � //$/6/H/Z/l/ ~/=�/�/�/�/�/�/ ? ?2?D?V?h?z?9 �?]�?��?�?
OO .O@OROdOvO�O�O�O �O�O�/�O__*_<_ N_`_r_�_�_�_�_�_ �?�_�?o#o�OJo\o no�o�o�o�o�o�o�o �o"�OFXj| �������� ��_'ooK�u�7o�� ����ҏ�����,� >�P�b�t�3������ Ο�����(�:�L� ^�p�/�y�S���ǯ�� � ��$�6�H�Z�l� ~�������ƿ����� � �2�D�V�h�zό� �ϰ��ρ�������� ۯ@�R�d�v߈ߚ߬� ����������׿<� N�`�r������� ������&�����	� k�-ߒ����������� ��"4FXj)� ������� 0BTfx7�I� [�����//,/ >/P/b/t/�/�/�/�/ {�/�/??(?:?L? ^?p?�?�?�?�?�?� �?�O�6OHOZOlO ~O�O�O�O�O�O�O�O _ _1OD_V_h_z_�_ �_�_�_�_�_�_
oo �?=o�?ao#O�o�o�o �o�o�o�o*< N`r1_���� ����&�8�J�\� n�-o��Qo��uow�� ���"�4�F�X�j�|� ������ğ����� �0�B�T�f�x����� �����ᯣ���۟ >�P�b�t��������� ο����՟:�L� ^�pςϔϦϸ����� �� ��ѯ���?�i� +��ߢߴ��������� � �2�D�V�h�'ό� �����������
�� .�@�R�d�#�m�Gߑ� ��}�����*< N`r����y� ��&8J\ n����u����� ��/��4/F/X/j/|/ �/�/�/�/�/�/�/? �0?B?T?f?x?�?�? �?�?�?�?�?OO� ��_O!/�O�O�O�O �O�O�O__(_:_L_ ^_?�_�_�_�_�_�_ �_ oo$o6oHoZolo +O=OOO�osO�o�o�o  2DVhz� ��o_���
�� .�@�R�d�v������� ��}oߏ�o��o*�<� N�`�r���������̟ ޟ���%�8�J�\� n���������ȯگ� ���Ϗ1��U��|� ������Ŀֿ���� �0�B�T�f�%��Ϝ� ������������,� >�P�b�!���E���i� k�������(�:�L� ^�p�����w��� �� ��$�6�H�Z�l� ~�������s������� ��2DVhz� ������
�� .@Rdv��� ����/���� 3/]/�/�/�/�/�/ �/�/??&?8?J?\? �?�?�?�?�?�?�? �?O"O4OFOXO/a/ ;/�O�Oq/�O�O�O_ _0_B_T_f_x_�_�_ �_m?�_�_�_oo,o >oPoboto�o�o�oiO {O�O�O�O(:L ^p������ � ��_$�6�H�Z�l� ~�������Ə؏��� ��o�o�oS�z��� ����ԟ���
�� .�@�R��v������� ��Я�����*�<� N�`��1�C���g�̿ ޿���&�8�J�\� nπϒϤ�c������� ���"�4�F�X�j�|� �ߠ߲�q��ߕ��߹� �0�B�T�f�x��� ������������,� >�P�b�t��������� ��������%��I �p������ � $6HZ� ~������� / /2/D/V/w/9 �/]_/�/�/�/
?? .?@?R?d?v?�?�?�? k�?�?�?OO*O<O NO`OrO�O�O�Og/�O �/�O�O�?&_8_J_\_ n_�_�_�_�_�_�_�_ �_�?"o4oFoXojo|o �o�o�o�o�o�o�o�O _�O'Q_x�� �������,� >�P�ot��������� Ώ�����(�:�L� U/y���eʟܟ � ��$�6�H�Z�l� ~�����a�Ưد��� � �2�D�V�h�z��� ��]�o���������� .�@�R�d�vψϚϬ� �������ϳ��*�<� N�`�r߄ߖߨߺ��� �������ӿ�G�	� n����������� ���"�4�F��j�|� �������������� 0BT�%�7� [�����, >Pbt��W�� ���//(/:/L/ ^/p/�/�/�/e�/� �/�?$?6?H?Z?l? ~?�?�?�?�?�?�?�? ? O2ODOVOhOzO�O �O�O�O�O�O�O�/_ �/=_�/d_v_�_�_�_ �_�_�_�_oo*o<o NoOro�o�o�o�o�o �o�o&8J	_ k-_�Q_S��� ��"�4�F�X�j�|� ����_oď֏���� �0�B�T�f�x����� [���󟷏�,� >�P�b�t��������� ί�򯱏�(�:�L� ^�p���������ʿܿ ���џ�E��l� ~ϐϢϴ��������� � �2�D��h�zߌ� �߰���������
�� .�@���I�#�m��Y� ����������*�<� N�`�r�����Uߺ��� ����&8J\ n��Q�c�u��� ��"4FXj| ��������/ /0/B/T/f/x/�/�/ �/�/�/�/�/��� ;?�b?t?�?�?�?�? �?�?�?OO(O:O� ^OpO�O�O�O�O�O�O �O __$_6_H_?? +?�_O?�_�_�_�_�_ o o2oDoVohozo�o KO�o�o�o�o�o
 .@Rdv��Y_ �}_��_��*�<� N�`�r���������̏ ޏ����&�8�J�\� n���������ȟڟ� ���1��X�j�|� ������į֯���� �0�B��f�x����� ����ҿ�����,� >���_�!���E�Gϼ� ��������(�:�L� ^�p߂ߔ�S������� �� ��$�6�H�Z�l� ~��Oϱ�s������ � �2�D�V�h�z��� ������������
 .@Rdv��� ���������9 ��`r����� ��//&/8/��\/ n/�/�/�/�/�/�/�/ �/?"?4?�=a? �?M�?�?�?�?�?O O0OBOTOfOxO�OI/ �O�O�O�O�O__,_ >_P_b_t_�_E?W?i? {?�_�?oo(o:oLo ^opo�o�o�o�o�o�o �O $6HZl ~�������_ �_�_/��_V�h�z��� ����ԏ���
�� .��oR�d�v������� ��П�����*�<� �����C�����̯ ޯ���&�8�J�\� n���?�����ȿڿ� ���"�4�F�X�j�|� ��M���q��ϕ���� �0�B�T�f�xߊߜ� ������������,� >�P�b�t����� ��������%���L� ^�p������������� �� $6��Zl ~�������  2��S�w9� ;�����
// ./@/R/d/v/�/G�/ �/�/�/�/??*?<? N?`?r?�?C�?g�? �?�/OO&O8OJO\O nO�O�O�O�O�O�O�/ �O_"_4_F_X_j_|_ �_�_�_�_�_�?�?�? o-o�?Tofoxo�o�o �o�o�o�o�o, �OPbt���� �����(��_1o oU��Ao����ʏ܏ � ��$�6�H�Z�l� ~�=����Ɵ؟��� � �2�D�V�h�z�9� K�]�o�ѯ����
�� .�@�R�d�v������� ��п������*�<� N�`�rτϖϨϺ��� �ϝ�����#��J�\� n߀ߒߤ߶������� ���"��F�X�j�|� ������������� �0�����u�7ߜ� ����������, >Pbt3��� ���(:L ^p�A��e���� � //$/6/H/Z/l/ ~/�/�/�/�/�/��/ ? ?2?D?V?h?z?�? �?�?�?�?��?�O �@OROdOvO�O�O�O �O�O�O�O__*_�/ N_`_r_�_�_�_�_�_ �_�_oo&o�?Go	O ko-O/o�o�o�o�o�o �o"4FXj| ;_������� �0�B�T�f�x�7o�� [o��Ϗ�����,� >�P�b�t��������� Ο����(�:�L� ^�p���������ʯ�� ӏ����!��H�Z�l� ~�������ƿؿ��� � �ߟD�V�h�zό� �ϰ���������
�� ۯ%���I�s�5��߬� ����������*�<� N�`�r�1ϖ����� ������&�8�J�\� n�-�?�Q�c������� ��"4FXj| �������� 0BTfx�� ���������/�� >/P/b/t/�/�/�/�/ �/�/�/??�:?L? ^?p?�?�?�?�?�?�? �? OO$O��/iO +/�O�O�O�O�O�O�O _ _2_D_V_h_'?y_ �_�_�_�_�_�_
oo .o@oRodovo5O�oYO �o}O�o�o*< N`r����� �o���&�8�J�\� n���������ȏ�o� �o��o4�F�X�j�|� ������ğ֟���� ��B�T�f�x����� ����ү�����ُ ;���_�!�#������� ο����(�:�L� ^�p�/��Ϧϸ����� �� ��$�6�H�Z�l� +���O����߇����� � �2�D�V�h�z�� ����������
�� .�@�R�d�v������� ��}��ߡ�����< N`r����� ����8J\ n������� �/����=/g/) �/�/�/�/�/�/�/? ?0?B?T?f?%�?�? �?�?�?�?�?OO,O >OPObO!/3/E/W/�O {/�O�O__(_:_L_ ^_p_�_�_�_�_w?�_ �_ oo$o6oHoZolo ~o�o�o�o�o�O�O�O �O2DVhz� ������
��_ .�@�R�d�v������� ��Џ�����o�o �o]���������̟ ޟ���&�8�J�\� �m�������ȯگ� ���"�4�F�X�j�)� ��M���q�ֿ���� �0�B�T�f�xϊϜ� ����ѿ������,� >�P�b�t߆ߘߪ߼� {��ߟ��ÿ(�:�L� ^�p��������� �� ����6�H�Z�l� ~��������������� ��/��S�� ������
 .@Rd#���� ����//*/</ N/`/�/C�/�/{ �/�/??&?8?J?\? n?�?�?�?�?u�?�? �?O"O4OFOXOjO|O �O�O�Oq/�/�/�O	_ �/0_B_T_f_x_�_�_ �_�_�_�_�_o�?,o >oPoboto�o�o�o�o �o�o�o�O_�O1 [_������ � ��$�6�H�Z�o ~�������Ə؏��� � �2�D�V�'9 K��oԟ���
�� .�@�R�d�v������� k�Я�����*�<� N�`�r���������y� ��������&�8�J�\� nπϒϤ϶������� �Ͻ�"�4�F�X�j�|� �ߠ߲���������� ˿ݿ�Q��x��� ������������,� >�P��a��������� ������(:L ^�A�e��� � $6HZl ~������� / /2/D/V/h/z/�/ �/�/o�/��/�? .?@?R?d?v?�?�?�? �?�?�?�?O�*O<O NO`OrO�O�O�O�O�O �O�O_�/#_�/G_	? _�_�_�_�_�_�_�_ �_o"o4oFoXoO|o �o�o�o�o�o�o�o 0BT_u7_� �oo�����,� >�P�b�t�������io Ώ�����(�:�L� ^�p�������e�� ӟ���$�6�H�Z�l� ~�������Ưد��� �� �2�D�V�h�z��� ����¿Կ������ ۟%�O��vψϚϬ� ����������*�<� N��r߄ߖߨߺ��� ������&�8�J�	� �-�?ϡ�c������� ���"�4�F�X�j�|� ����_��������� 0BTfx����m������$�FMR2_GRP� 1Z��� �C4 w B��	 ���;M8E�� �F@ c�5W�o�
8J��NJ�k�I'PKH�u��IP�sF�!��{?�  ���89�<9��896�C'6<,5���{A�  l/+BH5B�1�0 !@�33;"�33�7]/n-8/@UUT�*@9 � �{��>u.�>*���<���{>����>��l=�<��=�U�=�v!>1
{�:�ܜ:2B�8'Ŭ9IR�7���9f�� �/$?o/!?Z?E?~?i?��?��_CFG {[T �?��? OO�;NO �
F0HA �M@�<RM_CHK?TYP  ��p&(� ROMc@�_MINi@������@�T XSS�B�3\� 9�O���C�O��O�5TP_DEF+_Oz��&	W�IRCOMh@_��$GENOVRD�_DO�F��G]T[HR�F ddUdMTo_ENB9_ MP�RAVC]�G�@ �[F@� G��@GAw�\H͊#Iv0�Iά �?�Oo�o(oK* �V�QOUcPAqKRK<�@���oIo�o�o�o��C�  D�o�h1:A|A$ B�L.rpN�i�O�PSMT�d�Y*�@t�$HoOSTC�21eη@���7 M5C��T{���  27.02�=1�  e�_� q�������M�Ə؏���������	ano?nymous#�Q� c�u��������6�������F�'�9� K�]�o���������ɯ 쟆�0��#�5�G�Y� k�����ҟ���׿� ����1����g�y� �ϝ����������	� �-�p��ϔ����ߺ� ܿ���������H�)� ;�M�_�q�����Ϲ� �������D�V�h�z� |�R��ߑ��������� ���!3Eh��� �������*� <�N�PA��ew� �������// <n3/a/s/�/�/�/ ���/$/?X9? K?]?o?�?��?�?�? �?�/�?B/#O5OGOYO kO}O�/�/�/�O�?�O ,?__1_C_�?g_y_ �_�_�_�OT_O�_	o�o-o?o�~�qENT� 1f�y�  sP!�_�o  �p~o�o�o�o�o�o '�o3\�D� h������� G�
�k�.���R���v� ��鏬��Џ1��U� �N���z���r�ӟ�� �����ޟ,�Q��u� 8���\�����ᯤ�����گ;���_�"�QUICC0l�H�Z���~�1�������~��2����[�!ROUTER\�8�J����!PCJOG��χ�!192�.168.0.1�0��z�CAMPRYT����!��1��#�
�RTu�'�9ߚ�� !Softw�are Oper�ator Pan�elw�����`dNA�ME !mj!�ROBO���S_�CFG 1emi� �Au�to-start{ed�DFTP�O���O�_���O���� ����c_>�P�b�t� ���+��������� �@\�n��a���� x������ '9Kn���� ����O�O�O�OV ,/�k/}/�/�/�/v �/�/�/??B/�/U? g?y?�?�?�?�// (/*?O^/?OQOcOuO �OJ?�O�O�O�O�OO �O)_;_M___q_�_�? �?�?�_�O�_2Oo%o 7oIo[o_o�o�o�o �_�olo�o!3E W�_�_�_��o�o �����oA�S�e� w����.���я��� ��\n��s��� �����͟ߟ񟴏� '�9�K�]�������� ��ɯۯ�0�B�T�f� h�Y���}�������ſ �������1�T�ֿ�g�yϋϝϯ�����_?ERR g������PDUSIZ � V�^t�����>	�WRD ?�J�7��  ?guestV�I��[�m�ߑߣ���SC�DMNGRP 2�hJ�����7�V�8V�K�� �	P01.03� 8�   �e�?��  �;  �  �� ���������@�-��������x����0���y�d���`�,�>�P����?�  D���d����������_GWROU��i���Х��	���5{�QKUP�3�����V��TYC �����TTP_AUTH� 1j�� <!�iPendan��%`Ϗ�!KAREL:*%.@KCUew�M VISION SET����V�K��J( @:�^p������CTRL k�����%V�
<�?FFF9E3�5��FRS:DEF�AULT3,F�ANUC Web Server3* ! 5���1�C���/�/��/�/�/?��WR_�CONFIG �l�� 3/��I�DL_CPU_P5CR V�B�8�u0w BH[5MINf<�!�y5GNR_IO����V���]0NPT_SIM_DO�6��;STAL_S�CRN�6 ���I�NTPMODNT�OL�7�;�!RTY��8u1�6� ��ENB��7��Y4OLNK 1m��E�}O�O��O�O�O�O�OaBMA�STE�0��aBSL?AVE n��U�RAMCACHE�_�2O��O_CF1GI_`CaSUO��l_~]RCMT_OPR 8�2�ʟSYCLH_{U�L _ASG 1o��#�
 �Oo o 2oDoVohozo�o�o�o��o�o�o�o�K�RNU�M���
]RIP�F_XWRTRY_C�N�_{U�1���|A�b�� ]R�PfRp'^�=з=�]0P_ME�MBERS 2q���� $�%�r�����w��]0RC�A_ACC 2r���  V�Y� _ � �0� 5,P 6�JV�)��S�d� c�nU�  � 5��BUF001 2�s��= 	�u0  u0	�քU�ք�ք�ք�ք��փ

��+��;�L�[�m��|���������������Vփ~�~�!~�U1~�B~�Q~�c~��r~��u0( M��u0�`�x�u0I�+ט�~��~��u0�s8ր�uփ,���Cu0$Q�Yu04�@��d=��=PbVփq&��&��&�U�&��&��&��&�U�&��քքքU&ք5քFքVք�gքvք�փ��2 ��҃ց܁���� ��������ց� �����%��-� �5��=��E��M� �U��]��e��m� �u��}�ց������ ���������������� ����������Ő��͐ ��Ր��ݐ��吉�� ց������������ �������$�ց,� 1�5�1�=�1�E�1�M� 1�U�1�]�1�e�1�m� �u��}�ᢅ�ᢍ� ᢕ�ᢝ�ᢥ�᢭�ᢵ�ց��3ɯ҅� ��������� �"�#�"%�3�" 5�C�"E�S�"U�c� "e�s�"u���&� ���ҕ����ҥ����� ��ó��Ő��͐��Ր ��ݒ볢��&���� ��������� +�2�-�;�2�=�K�2� M�[�2�]�k�r�m�{� U�}���U򍢛�U򝢀��U򭢻�Y48�gQ2Et��4,%&�&��<&�K���25�H�IS��v�� ��S� 2023-�07-19Y& %|B;��p:�o� ����������������^W(V�sE�8Q� J\n���W'��Y!׀������s!�^��s  77��q5" 4FXj|��� ���//0/B/ T/f/x/�/�/���/ �/�/??,?>?P?b? t?�/�/�?�?�?�?�? OO(O:OLO�?�?�? �O�O�O�O�O�O __ $_~#�Ƞ/�A�S�b� dU��d3_�_�_ �_�_�_�_o!o! 3io{o�o�o�o�o�� c� �_��b� �-  L� 8  ^iO{OASe w������eO ,�+�=�O�a�s��� ��������ȏ�� '�9�K�]�o�����ʏ ܏�۟����#�5� G�Y�k�}���Ɵ��ů ׯ�����1�C�U�����T_f_S�"� X�Ŀֿ����� 0�B�T�BoTo�ϜϮ� �������ϿQ��� �Q��Q�� ������ f�xߊߜ߮������� ���?�Q�>�P�b�t� ����������)� ��(�:�L�^�p����� �������� $ 6HZl~���� ����� 2D�VhzCVI_CF�G 2wz� H�
Cycle �Time�Bu{sy�Idl�^�min}��Up��R�ead�DoYw�� ���Count�	N'um ����`,�w�7!EQPROG��xz���� p/�/�/�/�/�/?��@USDT_ISO_LC  z��p�J23_DS�P_ENB  �B;�c0INC �ys=w�P0A   �?�  =����<#�
O1�9:�o �1�?�?w��?�O\7OB� Cl3���6"AG_GRO�UP 1zB;�b<� �3�	nO�O?��/�Ow�Q �O�O�O_�O0_B_T_�f_��?IG_I?N_AUTO/D�:>c0POSRE*O<F�KANJI_MA�SK�V�ZKARELMON {z�h/w�y+_DoVohozoP�o�b�#|�'~3�w��e�_4KCL;_L�PNUMp0�o�$KEYLOGG'ING�`��bA{5�� LANGUAG�E z�Jp��DEFAUL�T Xqh�LG�Y}�*��w�x�0�  v�H [ �w�'0��w��w�?)7;���
�q(UT1:\�o� ��� �0�=�O�a�x��������(3o�c�LN_DISP ~�?���O�O��OCTOL9�w�Dz� K1�1>O�GBOOKq0i}�d���������X �|����ϟ����0us�'��	m��y�jA%;o�?�1k�_B�UFF 2�B; �w�2����� *2ү�� �-�$�6� c�Z�l�������Ͽƿ ؿ���)� �2�_π3~��DCS ��) �2�1$�c������������v�IO 2���� �3�jA�6�F�X�j�~ߎߠ� ������������0� B�V�f�x������������ER_ITM?>d�_?�Q�c�u� �������������� );M_q��8�I��SEV�`s=]�TYP?>.��!3��QRST�t�SCRN_F�L 2��� � �ϧ����//FDTPp??�C�NGNAMl4��Jrnr�UPS�GI\��U{5�!_LO{AD'@G %@*?%DMAYɥ�/�G�MAXUALR�M�b�QC��{5
��"�!_PR�$�P ha�%�� C��i��ٯè)3H@P 2]�w� �Ʀ	O!+t�0��0�P?�� �2�?�?�?�?���?+O OOO2ODO�OpO�O�O �O�O�O_�O'_
__ ]_H_�_l_�_�_�_�_ �_�_�_�_5o oYoDo }o�oro�o�o�o�o�o �o1UgJ� v�����	�� -�?�"�c�N���j�|� �����̏����;� &�_�B�T����������ݟ�ҟ���7��'D�BGDEF ��25?1>1@�R�_LDXDISAm ?+�MEMO_APg �E ?@+
 d����ү������,�>�� FRQ_�CFG �276h�A �@���!�<?4d%A���R�d��z2�2;�4�*��/�� **:�!���ȟ�!� ,�>�k�b�tϡϘϪ� ��#�25 �����'�� �6�,(��~���l� �ߐ��ߴ������'� �K�]�D��h���������*ISC 1�@)� �)�#��4 i�9�$�r�]��������_MSTR �����SCD 1��������,P ;t_q���� ��&L7p [������ /�6/!/Z/E/~/i/ �/�/�/�/�/�/�/ ? ?D?/?A?z?e?�?�? �?�?�?�?�?OO@O +OdOOO�OsO�O�O�O �O�O_�O*__N_9_ ^_�_o_�_�_�_�_�_��_o��MKg�������&o$MLTA[RMf��۷Qb �b��o�dQ��METPU��b�����NDSP_ADCOL�ef��noCMNT�o �e�FN�`�o�gFST�LIw�� ����g~�c���t�eP�OSCF5w�nPgRPM�o�yST�`�1��� 4��#�
����!�� !�#�5�w�Y�k����� ���ŏ׏����O��1�C���o��aSIN�G_CHK  �$MODAe���OkQn��DEV� 	��	MC}:�HSIZE���`ȿ�TASK �%��%$123456789 `��r���TRIG 1��� lQ�����`Lٮ��L�B�YP-��L�Ք��EM_I�NF 1�ۻ�`)AT&FVg0E0��k�)S��E0V1&A3&�B1&D2&S0�&C1S0=Z�)�ATZk�����H@ÿ�z�߯Ϣ�A�@C���g�Nϋϝ� Q� ��u��������Ͽ@� w�d�v�)Ϛ�U߾��� ���ߧϹ�*������ r�}�7ߨ������� ���&��J�\��� 3�E�W�i�������5� 4��X|�u �e�w��������0 B��f��EO� {��//�>/� '�/K�/�// �/�?�/'?L?3?p?��NITORPpG� ?�   	?EXEC1c�2U2�83�84�85�8T���67�88�89c�2:"D�2D�2D �2D�2D�2D�2D@ BDBDBC2%HU21H2=H2IH2UHU2aH2mH2yH2�HU2�H3%H31H3�2���R_GRP_S�V 1�@� (�w���<� ���>%��6�����u=���J�_D20�yS�ION_DBɐ�|͝a  �`fp O放T��`-��W�`Y`�!��qf0N   7�Z�P��[ pp�-ud1�/oAo�So�aPL_NAM�E !Q�|`��!Defaul�t Person�ality (from FD)�P��bRR27Q 1��L�XL�x<|a�P dzr�o �o�o�o#5GY k}������@���1�C���2�o n���������ȏڏ������<]�:�L�^� p���������ʟܟ�H �[i*�)�:�
)�^�]dPM��������� ү�����,�>�P� b�t�����g�y�ο� ���(�:�L�^�p� �ϔϦϸ����ϫ��� �$�6�H�Z�l�~ߐ� �ߴ���������� ��2� F@ G&h G��]gSP  �_�q�]bd[�C��������� D�7�Zj��	���=�@� -�X�N�`� r���������SP�0��4	]b-�	`B�<�N`:�oA�b���� Ag�  �	W�V]`-�S ]`��PC�T��s  h���)  �  u$�T&"�C �gyd���\k�R6R 1�ti�P�*0 � �f2|`  @D� � !?�#X�,?]`!]aA/���%]d.]d;�	�l,"	 �߀pJn ��NP`e  � � w� �� � ��"�SPK�K ���K=*�J����J���J9�٧�U�p��/SP@�_f��"j�@��(E14!�/�#�N����;f,1��� �a�������-�@¾ - T1�HZ0Z0� ��/  >c�=���>�]a���o���l? �?��2-!�3�&. Up�Pm P� ��P_�  ��P�F��*O�%	'� �� HBI� ��  ���&:��ÈlOÈ=�s�̈́E�"@�O@�@�>!�O/K"���&&�&�Q_  '�.T�!-0@2��O@����"=0@A?�C� C�PC��� Ca0Ce0Ci=�%��A�% 0� `l�-_hhX�'B�P��Q���A�U]aDz �on?3ooCoio�O��dIA�R�TZ��A����  �4@?��ff���o�ono  #{�!8�@9GzC>L�@�0(!�*(�@ uu�0�v�i{!t#t$�C�?]t�@,��<
6�b<߈;܍��<�ê<���<�^¬/�C�A�K"�#,"� �?fff?�@?&�&���@�.8���J<?�\�D�N\��I�R!�-$�)% |�'��
�`$�oЏ�� �ߏ��<�'�`�r�0]����He�F+P�� ҟ����m�����J���F�  F��~�BG�d GC�q V���R���ů���ԯ ���1��U�@��O�� �F�IG/�ӿ1���m� �0�B�T�:��o�{�33ϩ���ϸ������{An� ��_��EC��U��ϲ�d�?�؃ߊ��߮��Im�i4����C �CfPa0�¸�Ԑ0ؼ��@�@I���B�>�)A�C�A�IA��@?�?\����ú@ �������=q��A��Ay�I33@�0��@��C��1������(���C�����b��=q�Ů�����H��� G�� G��B�I��(E�ψ C�e�� I"�L�J�H�V@G5� E��x C��I3��J0�G��߀I�� 0 C ='�߀�k��������� ������"F1j Ug������ �0B-fQ� u�����/� ,//P/;/t/_/�/�/ �/�/�/�/�/??:? %?7?p?[?�??�?�? �?�? OO�?6O!OZO EO~OiO�O�O�O�O�O �O�O __D_/_h_z_�e_�_�_�_�_�_y�(΄�����r��<$e�U��o&o9�3�8�@oRo9я4Mgulo~o9Ѵ�VwQ�o�o4p�+4�]�m�i@�o(L:|u�P�r	P~~������_�0����{R��`G�2�W�}�h�  �`��ˏ���ڏ�����F�4�j�X� p�z��������ԟz����4�"�X�F�|����  2 F�@9�G&h�����9�B�&��)��C	�&�9�@-��9�o`�+�=�O��� ��{�Ħ�GAw\]�0����ɿ7�?��|p*9�t�9�9��9�{�
 ֿ9� K�]�oρϓϥϷ��π�������#�z�����hk�y��$�MR_CABLE� 2�hx i�ћqT�p@��¦�?>𦡆т����кƠ��C��ޱO�8�tB�����)ğ�+ޱFM�P��޴�ߕ��>��šz��C�N�|���=��a;�ް'E�mf�e����L�  ���C֠:��������a�_'�;bE��$T"�4��ՠ�y�ByМԡ��HE���ls=`޵;|�Vv�/� ����k������C�� L�>�8�f�\�n����� ��������?��H�� oq<���ܸ����ܸ*�,** \�OM ��i������޲^��%% 2�34567890	1i{ f��ް��ް�ްޱ�
�not �sent 5��WpuTESTFECSALG#�egۺ�d.$��Y
>$���p޴��޷Y/k/}/�/ 9�UD1:\ma�intenanc?es.xml�/�/�  ��D?EFAULTa�\ҿGRP 2�M � pė�޵  ��%1st m�echanical check�ޱ�z3鰄1�?��[ph��?�?�?�?��?޲R3controllerb4,O{?PO���?|O�O�O�O��OAMY=�O޲"�8SްQ_���kG8_J_\_n_�_�JC O�__�_�6/_o�o(o:oLoBC[0g�eW2. batt�eryPo�_�o��	 �_�o�o�o�o_i@�dui@ableN  D50Pqr�]�g�o������AddgreaYs;޷f��-ް�#���{P�b�t�h����A
ddoi�/��+�?��&�8�J�\�Adj7޶����<ް������
�؟���� �#|!too�����>ǟ��ய��ү�AOv�erhau�Ow��"� xް,�3�:5��`�r�������ްA$Q�пSV�� O� $�6�H�Z�lϻ���߿ �Ϲ������ �2� ��VߥϷ��Ϟ߰��� ����5ߝ��k��� d�v���������� 1��U�*�<�N�`�r� ������������ &8��\����� �������M" q�X�|��� ��7I/mB/ T/f/x/�/��/�/ �/3/??,?>?P?�/ t?�/�/�/�?�?�?�? OOe?:O�?�?�?�O �O�O�O�OO�O _OO �OsOH_Z_l_~_�_�O �_�__�_9_o o2o DoVo�_zo�_�_�o�_ �o�o�o
ko@�o �ov�o����� 1�Ug<��`�r� �������̏�-�� Q�&�8�J�\�n����� ��ȟ�����"� 4���X�����˟���� į֯���I��m�� ��f�x���������5��	 T¿��� *�4�F�X�j�|ώϠ� ������������0� B�T�f�xߊߜ߮��� ��������,�>�P��b�t����� � �b�?�  @�  ���	������H�Z�l��*��** @�>�7� ����������,>��e�^���A ���u���E Wi�Ugy�� ���/�/-/ ?/�/u/�/�/�� /�/�/??�/;?M?�_?�/�/���$�MR_HIST �2�>��0� 
� \
�$ 2345678901�?(�4�?���?9�)O ;O�?$O��O�O�O^O pO�O�O_�O�O_I_ [___6_�_�_l_�_ �_�_o�_3o�_Woio  o�oDo�o�ozo�o�o��oA�d�0SK�CFMAP  .>��08�1��`IYuONR�EL  �5�rq�0[rEXCFE�NB�w
psXu�qF�NC��tJOGO/VLIM�wd�3��[rKEY�w��_PAN�x+�'��[rRUN �,�SFSPDTYP�x<�uZsSIGN��t�T1MOT��q�[r_CE_GRP7 1�>�rs�2 ڰ9���c��8��8&� g����B�����x�� ��ڟ�ҟ?�Q��u� ,�����b�ϯ��ȯ� ��)�;�"�_�������|����7[qQZ_E�DIT��lw��TC�OM_CFG 1��h}�u�&�8� }
��_ARC_�r��5�yT_MN_oMODE����yUAP_CPL]���tNOCHECK� ?h{ @ ��������,� >�P�b�t߆ߘߪ߼�����ߍ{NO_WA�IT_L���ՀN�T���h{w��c�2�_ERR߁2�hy�1�6�����*���q�����w�O`�>g�| _ ���0�r�a<O�00 ?�5��O�5��p"�Y�PAR�AMa�h{���� ������1�� = O08Z lHx���������.��R~��ODRDSP\�����xOFFSET�_CAR�bψDsIS��S_Aw��ARK���OPE?N_FILE����;��S�OPTIO�N_IO!�3� M_PRG %hz�%$*E/W.�WO������p00�%�d.2  p��v� C�!	 ч�h�!�f����hRG_DSBL'  �7rqK�?�eRIENTTO��p�aC��pqqA� fUT_SIM�_D'or��hV~lLCT �<�粛$;��9�ed`7_�PEX���4RA-T� d�u�4��UP �q>��{ �OOOBOPI��$��2ރ�L��XL�x[3�0C�O�O�O�O�O �O__(_:_L_^_p_ �_�_�_�_�_�_�_ o�g2�O/oAoSoeowo �o�o�o�o�oB�o�o 1CUgy� ������f�o�~9@�!�N�P�K�]� o���������ɏۏ� ���#�5�G�Y�(�:� ������şן���� �1�C�U�g�y����� l�~�ӯ���	��-� ?�Q�c�u���������`Ͽ�s�¯��� � 2͠4A�!S�e�Gυ� ����A�����ϭ�������!�3�Q� W�uߗ���{ ��������	`����!�x�:�o@1?�Q�c�|u�A�  ��
V+��!+�21� �9���s  �h�p )  ?�  u$�� ���)��&�_�J����^fBl@O�01� �� � {D}��0 ��$�  �� @D�  ���?���X,q?+���+�D��������  ;�	�l��	 �߀pJ3 ������*  � � w� �I � �O�u�H(��H3k�7HSM5G�2�2G���GNɁ3h��(ϙ�u�C)H50�R50������r�û�¾  ��� �� �)���m�AK�µ�+�²���801 io���u����� p m�3�P00� �  � ��u��q�	'� � "�I� �  ����o�=���81/C+�@Y/_  Z�!�/��"������q�NA0�/  '�R0�$���CA0C�	��*C. ??�q��p�Az
b0�lwhhXn�B� �1��~�p!�5��zn��?3�?�?O .OU/GD!N2K4a+�Ӻ���@?��ff�ϏO�O3O !���O�KA8+��O�Z>LS ���J( +�:U�EV^I@99ң#?"T� ,A<
�6b<߈;����<�ê<�?��<�^�q�_2�AAp+���#���?fff?p ?y&�PD@�.�R�J<?�\�	bN\��U2�Q�@ ��Ao��`o�W%�O�o �o�o�o�o�o�o% 7"[mD�|��,oNoPo���xF��  F��+�G�d GCFQ�T�� d���u�����ҏ���� ����/M��&
 ������2�����d��J��O�[�3p ޟw�b�������
<�!A3�墚?+�C���x��w�)�?��H��O���s�
�4����C��C�࿇��b��b�a��@I��	B>�)A��C�AIA���@�?�\��������@ �������=q+�R!>�I�33@0��@���C�1����[�����C'��=q��Ů���	H�� G��� G�B�I��(E�� C�^l���I"L�J��HV@G5� E�x C����I3�J0��G���I�� E@� C��E� 0�i�Tߍߟߊ��߮� �������/��,�e� P��t�������� ���+��O�:�s�^� ��������������  9$]oZ�~ �������5  YD}h��� ����/
/C/./ g/R/d/�/�/�/�/�/ �/	?�/-???*?c?N?Ї?r?�?>�(I��ٙ^opR���5�5����?�?@�3��8�OO@�4Mg�u1OCO@��VwQ�]OoO4p�+4�]�M�I�O�O�O�O(_�L:�P�RPC^>�_�l_�?x_�_�_�_�[R�_�_o�_o,Bo-o  �@�EoWo �o{o�o�o�o_Q��o/{5?u c���?��������A�O�  �2 F@@�G�&hl���@�B�0���ձC��@�@򯷏ɏۏ����"�@��oL�^�p������@�?���AP@�J�d@�@�<���@�
 �����"� 4�F�X�j�|�������`į֯�?ʶ���-K��y��$PA�RAM_MENU� ?�E��  DEFPULSE���	WAITTM�OUTL�RCV�_� SHEL�L_WRK.$CUR_STYLJ�;��OPT�����PTB����C��R?_DECSNW�4U ���%�N�I�[�m� �ϑϣϵ����������&�!�SSREL_�ID  �E]Q��5�USE_PRO/G %0�%"߇�6�CCRc�G�]Q8����_HOST �!0�!���ߔ�T TP���ӿ�����4�>��_TIMEa�G����!�GDEBU�GE�0�6�GINP?_FLMSK]��qT�P���PGA��e |�;���CH��^��TYPE-�9�!��Q�z�u����� ��������
) RM_q���� ���*%7I rm������/��WORD ?�	0�
 	PyRy��SMAI����RSUͱ=#TE���S�	��J"CCOL�Uf)�/��LcЫ �@��`ȯ�d�q�TRACECToL 1��E:�� AP� ��'AP;P�.�&DT� Q��E0� �D � �� �[Q12��12�Ԑ12��12.5Ȑ10��]6_4_4	_4
�_4_4/2�54��=4�E4�M4�-4�*]6_4_4_4GЮ10� �4�4"�4�4���2_463�=4�E4�!`3.?@? R?d?v?�?�?�?�?�?��?�?E�D�A@��ED�MD�UD�]D���D�ED�MD�UD��]D�MVnC�}V~C���D��D��D��D���D�ED�MD�UD�J]D��D�}V�C��Du��D��D� 'T	'TU�O_#_5_ G_Y_k_}_�_�_�_�_ �_�_�_oo1oCoUo goyo�o�o�o�o�o�o@�o	-?�B�DU�D �D!�D"�D�#�D$?AN�  �O�O�O�O�O�OW	O O-K'1��o������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{�����k����� ����%7I[ m������ �!3EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_���_ oo1oCoUogoyo�o �o�o�o�o�o�o	 -?Qcu��� ������)�;� M�_�q���������ˏ ݏ���%�7�I�[� m��������ǟٟ� ���!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����� ����ѿ�����#���$PGTRACELEN  "��  ���!��7�_UP �����f��n�R�g�7�_C�FG �f�TP�!�g������ϸ�I���  ����{�DEFSP/D ��� �I���7�H_CON?FIG �f�N�W !�!�d-�M�F�  �0�P�����L�!��7�IN~~�TRL ��Ͳ��8��a�PE����f���,�\��7�LIDù���	��LLB 1��� �M�B�<�B4�� �M�%��Pպ� <o< �?�O� n�O�f������� ���"���<�j�P�r�����8������� 
Q�@3Ev�ٿGRP 1�����"�@��
����!�AM�D��@ D�@ C5f� @ �1���0�	�	,�,����uG���´F(BIpP:L�p��!�>�l7>�ú��/.� =�-=%�T/ Q//N/�/r/�/�/0/��/�/�/?)??  #DzN3W?!�
>?? .?�?�?�?�?�?�?�? !OOEO0OBO{OfO�O�O�O�J)�A
V�7.10beta�1�� A��=� R�!�A!��@�?!G�Q=y��#�B���$Q@�����B�l�4Q@�A���QT� �Oi_{_�_�_FTp���<��_�_�_�_ .� ��O��O�0oBo@,ofoPo�o�A-�p��u0�mf��o��o���@�AWP�R�c� B��B�>0uB�Hfs�d!�!�LPuM���d����r
�cx�tx��h��$|�����0��<�-�@�F�0�A��33`�������KNOW_M  ��"�����SV ��C�]�m? �� $��oH�3�E�~�!�����M��� �jR	��ѐlb���^���hhXd��1q� (�0u�8�4�����MR�� ���&�oj3�������OADBANFW�D����ST�1 k1�f��4�� �Y�!

��.�_�R� d�v��������п� '���]�<�Nϓ�r�@���ϨϺ����2��8��	�ݠ�<3�߂�3�/�A�S��4 p߂ߔߦ��5���������6�(�:�L��7i�{����8`���������MA֠���b�OVL/D  ��~��PARNUM � �������SC-Ha� o�
����8	�UPD�����#bb�_CMP_0��d����'�z�ER_CHK�����˒���RqSu�ٯ��_MO֯��_�a�_RES+_G����
V_�� ch������ �/
/;/./_/R/d/7�DT�/9o� �/�/�/;���/?? ;�!?@?E?;h�`? ?�?;���?�?�?;���?�?O;V 1���vߠ��@`}�\�THR_IN�Ru�f��dqFM�ASS~O Z�GM�N}O�CMON_QUEUE �����
�Qa�N U��N�F�H SEND8Q#YEXE._U�D BE-P_ SOP�TIOW,PPR�OGRAM %��J%P<O��RT�ASK_Ic�u^O?CFG ��O����_
`DATA���&kP�
2ʕyo �o�o�o�olo�o�o	 -�oQcu�:o�INFO���Wm� �DC����(�:� L�^�p���������ʏ ܏� ��$�6�H��w�t�Wl r)	a��K_a�i�~���ENBd�ѹ�2�ԘGa2̙�� X,		�=���� ���@�N�9�$��8�8�`D���_EDIT ��o����dWER�FLOXdC�RGA�DJ �}�A����?
���AϦQ�������??�  Bz��ga<8�
�v%$�\�è�r-�g�2���r	�H�@locBB=P���q@'�ǽ�*۰/ݲ *�*:�ֿ��q<��.@A��ſ�@K�@�c���\I)#����1�[ϩ�g�������w�A.@u����� ��O���K�5�/�A߻� e߷ߡߛ߭�'���#� ����=��y�s� �������������k� �g�Q�K�]������� ������C��?)# 5�Y���� ���1� mgy����� �_/	/[/E/?/Q/�/ u/�/�/�/�/7?�/3? ??)?�?M?�?�?�?�?{�	&o0OŠOWOBD�t$ qO�KEO�OAO�O�O	�PREOF ��ŠŠ�
ϥIORITY�W���ӡMPDSaP�Q��A�7WUT�V|��ΦODUCT�Q�}��O��OGg�_TG���R��vR�HIBIT_DO����[TOENT �1�}� (!?AF_INEaPo~g!tcpo>Gm!ud6oon?!icm^o��vRXY��}��š)� ��o�oŠ��o�e�o:! ^EW�{���@����6�H�*uS���A�J�����£�>Ԥ�Ѷ�/���z��¤�r�}�A~;�,  �P�}�8�J�\�n�ť�߆Zߏ����ҟ�£�]�ENHANCOE �i�}�A�AdޏD�+�rV�D� _�SɡӡPORT�_NUMbSŠ�.Uӡ_CART�RE���l	�SK�STAaW�[SLGmS`ٸk�;��HPUnothingL�)�;�M�]����������_�TEM�P څY���5�q�_a_seiban�OϯO(�N�9� r�]ϖρϺϥ����� �����8�#�\�G߀� kߐ߶ߡ��������� "��F�1�C�|�g�� ������������	� B�-�f�Q���u����� ��������,P ;`�q����������VER�SI@P�WQ �disable�^���SAVE �ۅZ	2670/H769'��!4���po� 	�	(kR�?;+2/ESe@O/x/�/�/�/�*g,���/z�n_�P 1ܸk�20
B�5�<?N?�7�@URGEb�B�P�^�aWFz0�QdT�pVW`�4LQ���WRUP_DE?LAY ݼ��5�R_HOT %�FnQ3�O�5R_NORMAL�8�R
O<_O.GSEMI>OdO|�O�AQSKIP3	�p�+3x�O_ _0_�M�5W_eWO_�_ �_�_o_�_�_�_oo 'o�_Ko9ooo�o�oYo �o�o�o�o�o�o5 #Ek}�U�� �����1��U��g�y��5�$RBT�IF�4��RCVT�MOUէå����DCR3��I� ��AC�}��C���C���?���>�9��<��Nä��`�`	1��$,��C`�	���OC�?_ <�
6b<߈;�܍�>u.�>*��<���U�p��?����� �� ߟ���'�9�K�]��o��������ERDI�O_TYPE  �!=����EDPR�OT_CFG e��G�4BH3�E���A2�� ���B� �T�b� ����:�����п��c� ϐO(�G_I�;�Y�[� mϣϑ��ϵ������ ߡ���E�3�i�Wߍ� {ߝߟ߱���	��-� /���?�e�S��w�� �����������+��� O�=�s�a��������� ���������K9 o]������� ��5#EGY �}�����/ �1//U/C/y/g/�/���/����INT� 2��9J��ǱG;� ?&;s���N?�f�0 l?~;�/ �?�/�?�?�?�?�?O O,ORO@OvOdO�O�O �O�O�O�O�O_*__ N_<_r_`_�_�_�_�_ �_�_�_o&ooJo8o no\o~o�o�o�o�o�o���EFPOS1 �1�̩  x�/:y�A?cN� �x-?y���� "��F��C�|���� ;�ď_��������� B�-�f����%���I� �������,�ǟP� b����I�����ίi� 򯍯����L��p� ���/���ʿe�w��� ���6�ѿZ���~�� {ϴ�O���s��ϗ� � 2������z�eߞ�9� ��]��߁�����@� ��d��߈��5�G�� �������*���N��� K������C���g��� ������J5n	 �-�Q��� �4�XjQ ���q��/� /T/�x//�/7/�/ �/m//�/??>?�/ b?�/�?!?�?�?W?�? {?O�?(O:O�?�?!O �OmO�OAO�OeO�O�O��O$_�Cu2 1� �O�O_�_{_�_�O �_s_�_�_�_2o�_Vo �_zoo�o9oKo]o�o �o�o�o@�od�o a�5�Y�}� ����`�K���� ��C�̏g�ɏ���&� ��J��n�	��-�g� ȟ��쟇����4�ϟ 1�j����)���M�֯ q�����ϯ0��T�� x����7���ҿm��� ��ϵ�>�ٿ���7� �σϼ�W���{�ߟ� �:���^��ς�ߦ� A�S�eߟ� ���$�� H���l��i��=��� a����������� h�S���'���K���o� ��
��.��R��v #5o���� �<�9r� 1�U�y��� 8/#/\/��//�/?/ �/�/u/�/�/"?�/F?<,_>T3 1�I_�/ ???�?�?�?�/O�? )O�?&O_O�?�OO�O BO�OfOxO�O�O%__ I_�Om__�_,_�_�_ b_�_�_o�_3o�_�_ �_,o�oxo�oLo�opo �o�o�o/�oS�ow �6HZ��� ��=��a��^��� 2���V�ߏz������ ��]�H������@� ɟd�Ɵ����#���G� �k���*�d�ů�� 鯄����1�̯.�g� ���&���J�ӿn��� ��̿-��Q��u�� ��4ϖ���j��ώ�� ��;�������4ߕ߀� ��T���x�����7� ��[������>�P� b������!���E��� i��f���:���^��� ��������eP �$�H�l� �+�O�sY?k44 1�v? 2l ��/2/�V/� S/�/'/�/K/�/o/�/ �/�/�/�/R?=?v?? �?5?�?Y?�?�?�?O �?<O�?`O�?OOYO �O�O�OyO_�O&_�O #_\_�O�__�_?_�_ c_u_�_�_"ooFo�_ joo�o)o�o�o_o�o �o�o0�o�o�o) �u�I�m�� �,��P��t���� 3�E�W����ݏ��� :�Տ^���[���/��� S�ܟw� ��������� Z�E�~����=�Ưa� ï���� ���D�߯h� ��'�a�¿��濁� 
ϥ�.�ɿ+�d����� #Ϭ�G���k�}Ϗ��� *��N���r�ߖ�1� ����g��ߋ���8� ������1��}��Q� ��u������4���X����|������5 1�M�_��� ;A�_����� T�x�%�� �j�>�b ���!/�E/�i/ /�/(/:/L/�/�/�/ ?�//?�/S?�/P?�? $?�?H?�?l?�?�?�? �?�?OO:OsOO�O2O �OVO�O�O�O_�O9_ �O]_�O
__V_�_�_ �_v_�_�_#o�_ oYo �_}oo�o<o�o`oro �o�o
C�og �&��\��	� �-����&���r� ��F�Ϗj�󏎏��)� ďM��q����0�B� T����ڟ���7�ҟ [���X���,���P�ٯ t�����������W�B� {����:�ÿ^����� ��ϸ�A�ܿe� �� $�^ϿϪ���~�ߢ� +���(�a��υ� ߩ��D��߳���6 1� ��zߌ���D�/�h�n� ��'��K�����
� ��.���R������K� ������k������� N��r�1� Ugy��8� \��}�Q� u��"/���/ |/g/�/;/�/_/�/�/ �/?�/B?�/f??�? %?7?I?�?�?�?O�? ,O�?PO�?MO�O!O�O EO�OiO�O�O�O�O�O L_7_p__�_/_�_S_ �_�_�_o�_6o�_Zo �_ooSo�o�o�oso �o�o �oV�oz �9�]o�� ��@��d����#� ����Y��}����*� ŏ׏�#���o���C� ̟g�🋟�&���J� �n�	���-�?�Q��� �ׯ���4�ϯX�� U���)���M�ֿq���<����7 1��ߧ� ���q�\ϕϛ���T� ��x���߮�7���[� ����,�>�x����� �ߘ�!��E���B�{� ��:���^����� ����A�,�e� ���$� ��H�����~���+ ��O����H�� �h���K �o
�.�Rd v�/�5/�Y/� }//z/�/N/�/r/�/ �/?�/�/�/?y?d? �?8?�?\?�?�?�?O �??O�?cO�?�O"O4O FO�O�O�O_�O)_�O M_�OJ_�__�_B_�_ f_�_�_�_�_�_Io4o moo�o,o�oPo�o�o �o�o3�oW�o P���p�� ���S��w���� 6���Z�l�~����� =�؏a����� ����� V�ߟz����'���8 1�*�ԟ� � ����¯ȟ毁�
��� �@�ۯd�����#��� G�Y�k�����*�ſ N��r��oϨ�C��� g��ϋ�߯������ n�Yߒ�-߶�Q���u� ����4���X���|� �)�;�u�������� ���B���?�x���� 7���[���������� >)b���!�E ��{�(�L ��E���e ��/�/H/�l/ /�/+/�/O/a/s/�/ ?�/2?�/V?�/z?? w?�?K?�?o?�?�?O �?�?�?OvOaO�O5O �OYO�O}O�O_�O<_ �O`_�O�__1_C_}_ �_�_o�_&o�_Jo�_ Go�oo�o?o�oco�o �o�o�o�oF1j �)�M������0��T�:�L�MA_SK 1�W�N������x�XNO � ������MOTwE  ǌ  ��_CFG ���O�l�PL_RA�NG ��q[��A�O�WER �W��y�`�SM_DRY�PRG %W���%����TART� �q���UME_PRO�����H��_EXEC_EN�B  �t\�G�SPD��6�>��K�TDBY�k�RM�z�k�IA_OPTgIONQ��^���INGVERS���Ȋ
�o�I_AIRPURO�� ��Մ1�m�MT�_��Tl��`�OB�OT_ISOLC�Ō�-�4�0�o�N�AME���n�OB_CATEGň�y�փ̀���سO�RD_NUM ?�q�*�H?769  �t@��R�d�x�PC_TI�MEOUTQ� x�x�S232�1��ȅj� LT�EACH PEN�DAN���8����Ƽ ��pMa�intenanc�e Cons�r�����"���tNo Use�����@��R�d�v߈�v���NPQOΐ��8�̥��oCH_L���^��J�	���!U�D1:1���R�VgAIL!�¥�\���SR  ��ʡ8���R_INoTVAL���\���໮��V_DAT�A_GRP 2�|ȅ�� D��PL�/�H�S�>�ȅv� ��n������������� ����F4jX� |������ 0TBdfx� �����//*/ P/>/t/b/�/�/�/�/ �/�/�/??:?(?^? L?�?p?�?�?�?�?�?  O�?$OO4O6OHO~O lO�O�O�O�O�O�O�O� __D_́�$SA�F_DO_PUL�S���p[��SC�AN}���[���S�Cm�� �`�Xj��p�p
��1�`�(�վQ�r H��_ oo,o>oPo�_to�o`�o�o�o�o����Eib2�d�Q�Qdx��a
q�	�T�i @7�FXjtv&y:� ��t�_ @�sTʠ������T D�� �+�=�O�a�s����� ����͏ߏ���'��9�K��߯�8w�Z�����n�  ��;�o��ʑ���p����
�t���Di_�jaѰ�X � �����U �Q9�K�]�o������� ��ɯۯ����#�5� G�Y�k�}�������ſ ׿�����1�C�U� g�yϋϝϯ���������	ߗ���2�D�V� h�zߌߞ߰�����e �� ��$�6�H�Z�l� ~�����}�0�r� �&�������)�;� M�_�q����������� ����%7I[ m������ �!3EWi{ �������/ ///A/S/e/w/�ߛ/ �/�/�/�/�/??+? ������ibk?}?�?�? �?�?�?�?�?OO1O ?IROdOvO�O�O�O�O �O�O�O__*_<_N_ `_r_�_�_�_�_�_�_@�_oo&o8o,x�a� �Co�o�o�o�o�o�o �o�o"4FXj|���zmo��.�v��+�����	123456�78]2h!B�!��%�\1}�k`�T�f�x����� ����ҏ��lo�� 1�C�U�g�y������� ��ӟ���	��-�>� ��a�s���������ͯ ߯���'�9�K�]� o���@�R���ɿۿ� ���#�5�G�Y�k�}� �ϡϳ����ϖ���� �1�C�U�g�yߋߝ� ����������	��-� ��Q�c�u����� ��������)�;�M� _�q���B�������� ��%7I[m �������� !3EWi{� ������// //�S/e/w/�/�/�/ �/�/�/�/??+?=? O?a?s?�?McE��?��?I/�?�?O��Cz  BpIj �  �H2_b� } 6�F
[G�  	�AD�?�O�O�O�O�K	Do�<�uO_$_6_ H_Z_l_~_�_�_�_�_ �_�_�_o o2oDoVo ho�O�o�o�o�o�o�o �o
.@Rdv �������#���B�1iA�<�� �iA  �/�I��v,�mAmAt  6@m�����x`�$SCR_�GRP 1��*P30� �� ��A ��	 Ё�؂���1 ����w��#��J�Mg�K@G�DCv����N�G��L	�M-10iA/8�L 123456�7890k@�� �8k@MT20 L͐-C
ș��,�A^H �؁Z�@ǁ'�ǁ�C�G���-�	�v����������ά��H�؀_�܇ǂ���� 5�G���o�A"����������^� h�@,V�U  [��B�%@��������A6@ �  a@�@8��N�?�^����H%@q�K��F@ F�`�£Ϛ� �ϲ�������!��E� 0�i����8�h���ߣߵ�B���X�	� ��-��Q�<�N��r� ���������O�q�3�!�F��]@C�x�x�B`�8�>���~�D6�i�@8���%@���ȗ�'��?-DCA��1a�]�> �A2�A T{���
i���� (� � $ ��H3l)J��Γ���ECLVL��A���7�?A��*SYSTEM*�@�V9.10214� �8/21/2=0�A �@��z�SERVEN�T_T   $� $S_NAM�E !	 PO�RT�@!ROT�O! �_SPD�  ��/ T�RQ   
^,#AXIS5!:'�2  2c�,#DE�TAIL_ � l $DAT�ETI! ERR�_COD�#IMP�_VEL4@ 	�"TOQ�$ANGwLES�$DIS���&" G%%$LI�N�"��,#REC�5! ,!O%i � MRA�! 2w d2IDX�"��$B  �0$�OVER_LIM�I I 	+$OC�CUR5!  ��+COUNTE�R! + FZN_�CFG5! 4 $ENABL�#�ST� "FLAG^"DEBU�3R�!�� � �1��5! �� 
$MIN_�OVRD�@$I��� �2�1�5FAC�Ee"�1SAF�7MIXEDL�9�!�2�ROB%$NE�&APPx2�SHE�LL�4	 w5$J?@BAS�#�RSR_�5  ?$NUM_y@� � xA1�'y@2��J3�J4�J5�J6ʜJ7�J8�'lARO�O � CO�ON�LY�$USE�_AB#xBAC�KENB�  PIN�>0T_CHKSO?P_SEL_�0,Yg_PU;Qo1M_�!;OU#PNS|F P�YC�&�0EPM�%TPFWD_KAR�!� P�!RE$$O�PTION�2$QSUE�Y" D�RYRB�$CSTOPI_3AL;SYCEX+STQl�P�$XTSPM1i�2"MA�1STY�;TSO
`NBRDIGQTRI�3�Q�W�INI�M& 8bNsRQxf`ENDNd�$KEYSWI�TCH�S�QZa�TH}E�PBEATM�SPERM_LE�"R�QE� �gU�SFd��RS_dDO_HO�M�0ORA/PEFP0 !"0�3U ST�bR�C�`OM�#�!OV�_MSJQ ET_IOCMN+S�W5a��XEHK !
 gD �7qSU�"f�RMP+S� PO7B�$FORC�SWwARNQ��XE�OMrP 7��$FUNC��3UL	0}QAR'`�u2�vE3�v4�qorC0O�P�L�r�"�XUNLiOeP�$:�ED� ���SNPX_�AS�2 0�@A�DD�0�1$SI}Z�!$VAR�'�MULTIPR�Z��pA�q �� $tY[�r	��B`�"�AC� ΆF'RIF">0S�P�y�"t��NF{dODBUS_ADw2�B���&CM�aDIA��q$DUMMY�15aM�3J�4J���Sz@  � Lx��"TEqM�8J��SGL��TAJp  &�0���@J�<����STMT�Q���PSEGb��BW<�P��SHOW��!�BAN̐TPOF��M�9J�0J�(a�+ VC�G�2 ��$PCpP?0-�G3�$FB�qPD�SP"�PAFPF�)�D/��2�� ��!A0��@� ���p���p���	������5��6���7��8��9��A��B���p��h ��Ր��F���P���T�P�P��l�P�̩1٩1�U1�1 �1�1�U1'�14�1A�1N���!ǘ�2��2��2���2̩2٩2�2��2 �2�2�2�'�24�2A�2N�3���3��3��3��3���3̩3٩3�3��3 �3�3�3�'�34�3A�3N�4���4��4��4��4���4̩4٩4�4��4 �4�4�4�'�44�4A�4N�5���5��5��5��5���5̩5٩5�5��5 �5�5�5�'�54�5A�5N�6���6��6��6��6���6̩6٩6�6��6 �6�6�6�'�64�6A�6N�7���7��7��7��7���7̩7٩7��7��7 �7�7�7*'�74�7A�7N���VP�`U3" Q< �B
��V�� ! x $T�OR�Q@�  �"Mb$ R1 L@BQ_W0AR��%T!�p�$S[iC�Qp�_U�^��8��L� >  � x�� �7��m��0���`�R�VALU�5QP�V]z�F�ID_L��"%HI*I�r$F�ILE_xSM$BD�$sN0�SA21� h5y E_B�LCK�S�"���(D_CPU�)y��)m���3P/b$q�Y��rSR�  � PaWY0P�� 1LAƑ�S11314RUN_FLG(54,1�4�`/5M14M15H`rP4o04'�T2�Q�_LI�r  ]k@G_Ob�P�P_EDI+Rq�T2 @�3�20�$P��!����TBC2x� �}�8P/0T�Q�1FT'dD5cTDC/0A`a�0@aM	�F.AGTH�"��DDOPGRQH��pERVE(crD5c�rDa��14PG@ �X -$�AL�EN(c�D5c�@`R1A�PF��W_k�#i1�A:$2�GMO�!C�S�DPIZP�F!0Y8�@![DE1U��LACEXrfCC8B���`_MA^�0V8jU@WjQTCVq\�Q@WT�a�Z�U�Zd�/SP]��U@S]�J@`AG��M�T�Jjgv�/Ua@U�A2)pp\��5a.SH�JKHfVK@$�ZaU�Zaa�O`J�lra^cJJfcJJncAAL^c�`fc�`�fdm��b5OC�PN1�\P�`�[nP�L
P_���m!�0CFb� =`5GROU ����P�N�0C�� pR�EQUIR]B�E�BU̓�A�V$T1P2Vq�@@v�1a���4 \�p�8AP�PRLpCL�
$:�0N�xCLO�0�y�S:E�y/U
�1�� ��0M,@oP�PF�N�t_MGI��pCx��z �d�lP�BRK��NOLD��R�TMO�1I�6��uJ�0H�P�dLPfcLPnc�LP�cLP�cLP6��7ȃ����p�B�4G� Ir�B$��<U��PATH��@����H��p[p�.�SCA�2L��r�qIN�BUCP�A\�-Cf�UMe�Y�@� `l�&!xA�����������PAYLOA�D�J2LR_A	N$AȓL0ҙΑ�ޑ�R_F2LS3HRlD�LOӔ[���i��i�ACRL�_�!Y�L�U���gbH���$H�z�F�LEX�s�0J�6 P�r�?
OqO��Om"���E  :�O�F@P�#��Oha0@P�O�O�LF1#�q� ���O__0_B_T_��E^_p_�_�_�_�_�_ �_�_�ȩ��WcHd��@��o!o3o"�:jT����XraFe���Qe Z�3�]ooo�o�`�e�e@�e�e�o�o�o�j	��t! ��0#5�B@AT��Hq�PE�L�T1p�OxJ[p vVpJE3�CTRU�ƙ�TN)l�@wHA_ND_VB���� ׄ" $��F2��<D�SWl"���q�v#� $$M��yM#��2�-�O� �q�K�A) ���v�(!h� �A��#�A�1�A@�s��� #�D*1�D@�P �G"0		CST%�2�NC�DY.0�p�T�{��� �@�#�����Hg��K�-�G�P���������������ʂЂJ�5$c ���� Ʊx�qASYM0��Ip0�#wL��P�_n0A�a�t�^�`@��~�������ƓJ͜�~�ߚ������_V�I��<(�sM V_�UN�2; b#��
�J Iez"�z"�~$4��$ �&=��PP�~�_�q�5�;��������0HR�0�1%��01���2DI@�;sOO4�210N�& �Ђ�IeA��4�|1����3���|���20 ' �� ��ME����Х2�"�TC0PT@����1�`������8�1�9T��a� $DUMMY}1��$PS_���RF^��`$(Fn�pFLApYP2��BB�3$GLB_�T�E5]E�0��_�8ڱ��1( X�p@w�ׁST��VpSB}R�M21_VRrT$SV_ER�1O��C�CCLw@�BeA�O2,0GLD ;EWq) 4p�1W$Y��Z��WS>`���A�0e��r�A]U�E* ��N P��$GI��}=$�A )р�APq+ LpAV��}$F�EIVNE+AR�N��F�Y��TANC���8��JOGR�t� �,^0$JOIN�T=�N� �CMS�ETq-  >WE(vU�:�SA��[T;�q.� ��U���?�VpLOCK�_FO���K0BG�LV��GL:hTE�ST_XM�p�QEMP�PRr^buB%`�$U��B=�2*VpS�a+Ob��*`�a�)�ACE�`RS�` �$KARP�MQ3T�PDRA�@�d�QVcEC4��f�PIU�a�,�aHE,`TOOiLe��cVd�RE�`'IS3�r6�����ACH�P[p-qO�>��3D3��QPS�I�r  @$R�AIL_BOXEz=��@ROBOUd�?��AHOWWA�R��tq%@@qROLM0B�u �=t�r0�bp܍�ـO_F1�!>�@HTML5D1U�G�	c2qځ/�^� �R�`O��0��R]��Q�p0@�CO�U�R1 d�@�e)��v�P�%`$PIPVfN0�rbr2q����a�p�CORDEaD*`6���PXTV��DQ),0,�O�0 �2 D \@OB ��z�*`����C[@��ܶ|�SYS��ADqR{�,0�0TCH:�� 3 ,��ENT52��A1a_AT�x	���'�VWVA�1?4 � �`�B�E5PREV_RT~�$EDITT�_VSHWR1��F(s�� Q< D�0������$HEA�D�� ���\�K�E Q@CPSPD���JMP��LD5g�TR�g45��T���I_`S{�C���NEp|��TIC)Ke�oM���A�{HN�A6 @��8��Ñ_GPR�Yvγ�STY	�>qLO�wA(S�N� �7 tk 
O�G�%$4��AT=�@Sq�!$@p!=м1HEy0GFPRR�SQU�`X�IB;!�TERC�0Q8�{TS�8 HP��@.�0�-���a}�O�0�3��IZJDAQFE$APR��1Ap����.�PUAဵ_DO��R�XS�PKD6A�XI���s�aUR I��|�{p@�͆��J�Y_�`߂ET�P3b���5��F5��A,B8D9Hw���Up`2SR��9l ��M�%�[�8�m� K�[�V�[�d�[�t��� ���Ŧ��Ŷ������������!��C6���C��ͯ����qSS}C_@ : h�@cDS`��a@SPv0&��AT��L���?���BADDRESzsB_�SHIFA�^{`_2CH{�Ɂ�I~@��TU~@I�*� ;�RCUSSTO�&�VbIj2A< �Gh��d�
^j�
��V-����0= 	\�@G����o�>�����C��A��~�F��B����TXSCRE�E��><0��TICNA�COP��AT,�8���? T���@ d�߁�A�@L���ނ��H�[�RRO �Pހ���E�Ŵ��UE�@# �-��6@S�A߁'RSM?���U��
�D6��00S_S��i ������i�Cb���3� 2?*PUE�Ap2�Bp�GM�T� L�!���@O~�U �BBL_Bp9W�0�0B ���v5OQ�LE�xzpE�RIGH��BRD�D�CKG�R�0�T����WIDTHHs��ĲUq|BAq8�UI�pEY�Щ1C6��p�p�bpl�BACKЀ�0B1�A�0FO��DLAB��?(�0I@p#b$URL�qqCO	�0Hl� D 81�P_����0R P%b/ÔHx6��O�0E�I��G� U� �R3b�qLUM�Ķ�GERVM��@
P�PjF�0�GEu0{Q������LP4%
�	E���)Q'��_(�Ѩ_(,p^)5\+6\+7\+8A"��3k��P���F,qaS��E�	USR�DG �<�@�0UERT�ERF�OB�ERPRI�mxLp�!30TRIP^qm�UNDOg5H<PàL0���q����{bްؠ I��� o�G ��T0�p�� �2OS�1�6AR�r�v3�a�AJ�O@S^�2b���{bU<!�AK�?�?��<"a�v3�OFFT`�@L�@z�3OU@ 1J�@�?DgDK�@GUفP�fA��C}ьGSUqBb��@/ SRT�0�B�MI��Q�pO�OR�Bp�ERAUT��DT��I��A_R��N 9|]��OWNy0�$SRC}������DT`>UR�MPFI8y�y��ESP|�G� �u#��'r�BQ�m�6O `@WO���=��COP&!A$հ{0_YPrX�Q.��UWA_�Cra��Q�P�S�Qr ��4��rW� P?�SHADOW��s"a?_UNSCA�c"c��/cDGD7q��E�GAC�Sd��PP�G�Q���ST�E���O��t�P�E"��VWDt�F1TRG�6R y�>��jMOVE}�#A�bANG���f-C��f�3�bLIM_X !Cv'Cv�hq|��`�g?06��`"BVF�М�Cs1VCC���S?�C��RA���`ϥ\D��@NFA�R@�Z]�E,�Q>0G��f��R:�{0DE�b��p���p6T�# i�؁ϣ�u��㡹W C% �DRI�`��aV[�*���S�D�$MY_UBY�$�}�3ϥ~���b�����Q��P_8`�y���L��BM��$�DEY
�EXXc ���UMUِX�d�����US��˰.0_AR�"B#06��fG�PACIqt�`HQ�d�I�-CI��3I����QR!E���1f�sI�N�U ?�PG�`!P�⎐. �sR�0�AV�k���B	�R��R�dSWA�osh I��n�O�!�A��[�E� U���ah Y/��sHK��W����aS���Q��cE�ANS��P��+�MwRCV6X �- UO�pM�C��	��8?C����REFb�� ����
r�ِ0���@��꡹����A�_;P W�B�o����`��k�\����x�r`�r3Y ���a��ϒ�1`�$GROU���3��¶��s�pT����20$0 ����0X V�Ӂ�Xֱ���UL�qW�P�C%p�X��NT�S+ĔR*��6��!6���L��_Ű�_���k��!�pTIЙ�Z� t@MD�@AP�_HU�q�`��SA.Q�CMP}�F�����Ų�_��Rqty����W�j�X��F1VGF|`S[� �qM0����UF_{�0˂��@JʼRO� T��շ����|.�UR1E9��6�RI;���I&༨�o�o{FQyXFQ'C`wIN�H��xx� V�1,r��A��?�W�|��Q/��V����LOp'�\ax ������!NSIIBV�IA_�R;�\ ��� HDR )�$JO� b��$Z_UP)p��Z_LOW�������\(p���P鱬3�9���Ⴐ��'Q�| �"�]� 0��PA� �CACH���}���퀙��!�P]SC(qIB�F�#���T� ��|�$H	O�1R��/�%�" f������?�RQ0!���cPVP���pH_SIZ�sRZ��M��N�Q�MPr
�qIkMG�d��AD�	��RMRE���WG�PM�pNDRP�VA�SYNBUF�VV�RTD� W��OLE_2D,tc�J1@C�qUۃ��Q���ECCU{�VE�Me�}�d��VIR�C��
" {�L�A��RQ}0\0��AG:R�XYZ)��C�W�������A�T�p܂IM��|G`��GRABB�1�Y�b2b���^{�>
�CKLAS�¡8b�Y@_  񱵵IT��5P@�21T$b��p!�` ���SP�G�%TQ�RQ�q�P�"�x�I�$|��=�BG�_LEVE�QL�PaKL��"ѥ�GI� �NO�Q܁��͐HO|bPRa � �F����E6S��g]2{ROQ�ACCEe@���px4VR�A��y1܂R`� AR�cP�A@�>��D�SRE�M_BQ$�p�"JM�PU�XAbi$1�$SSlSFD�Ќ"����Y@c  ��S�� ��N/DS�VLEX�&dbSdqg`,��&DR�w$YQqH�(`qH҄�c ���VP2h�e�� �є`V��cPMV_PI��DX�`��@3����IF&�\rZ �JT�E�@���H���E�AGAU?�LOO�d?�JCBTZ�'Bx`H +cPLAN'r��L2��Fw��D?V5Y �WM��~Ppu�T�FS��U�Q�ѥU�� ��V2DbX�1L�RKEZq�1VAN9C]C�R_O�|`f (�p8�s$\��3Zr��R_A3� g 4��dovn#pp� �_���h h�p�9��ĬvOFF�safW@�����EA��Y
� LSK��MN��q�g S`��|@>c"i < WJ��^=�UMMYY����\�D�P�AC�U��1�U�pj �$�TITV1g$PR8A��OP�����SF���Cki ��|6����!SMO"!�l%BXC�4J�p�v��ZD�vm DQx6�AL^1IM; ���0IN�MSG_�Q�Sw
���_w�pn%B�w�8�%�M� �XVR�"�oI"�pT�5��ZABC���p��Ƃ��Ӡ
 �Ā&��`VS.� q � w0���=�CTIVeAI�O�b�	s�ITVlLW�DV@
l�"��2� DI�� @�� ��|A��d���N�LSTs���ݰ��7_ST��A%��DCSCH��r LQp�����~P1��m�W GN����r���_FUN�� �A7ZIP!�s%B� �L8�L|�Ѣ�aZ/MPCFʅt�r9����L�DMY_L�N$pq��M&�˄u $��Q��CMCM��CLCOART_����P�a? $J����D=��¢��u�ǥu����_�����U�X�P�UXEUL ����
�̥
��.�8�>���FTF����k���m�Z�vC �*����Y%��D.  w 8 �$R� U�Q��EgIGHe3�x?(�0Ԛ�0���P@%x a�=0�sq�$B������b_SHIYFB�	�RV�PF��&1�	$)0C�ঢ ���d�pl��r�"l���D|ȕ�C �NV:�a��SPH�0%чy ,�0��ֿ���$S{0DEFAU�n�B����������HOT䣐����MIPOWERFL �@�����%�WFDO�� ����Y��`?1 ���q��� L!ip_E�IP5ԑ����j!�AF���`�߼�!'FT�������3!��-����S�!R9MHQp�7灺B��f��po�5������!OPCU�A�����7�!�TPP�@8���d<&���!
PM�p�pXY����er���J�����f��!RKDM-@V��g
>g!R90h��hV�!
h�~�����i��!RL�SYNC &8|�K!ROS���r�4:�!
C�EL�MT�`���kL��!	��PS����l�//!�WOASRC6��m/v{/!�USB|/��nj/�/!STMP��/��o�/?�7?*?`=e�I��K�L ?%q� (�%SVCPRG1`?�:�52�?�?�03�?�?�04�?�?�05 O%O�06HOMO�07pOuO�08�O�O�0	9�O�K�4~�O�1 �?_�1�?=_�1�?e_ �1O�_�1:O�_�1bO �_�1�Oo�1�O-o�1 �OUo�1_}o�1+_�o �1S_�o�1{_�o�1�_ �1�_E�1�_m�1 o��1Co��1ko� �1�oe?w2�0~?�00� u��1y���������� Џ	��-�?�*�c�N� ��r�����ϟ���� �)��M�8�q�\��� ����˯���گ��� 7�"�I�m�X���|��� ��ٿĿ�����3�� W�B�{�fϟϊϱ��������k:_DEV �q��MC�:�4���GRP 2q����0�bx 	� 
 ,c��|�<� hߥߌ��߰������� #�
�G�Y�@�}�d�� ���������d�1� ��U�g�N���r����� ������	��?& cJ������ ���;M4q X������/ �%//I/0/B//� �/�/�/�/�/�/�/�/ 3??W?>?{?�?t?�? �?�?�?�?O�?/OAO �/eOO�O�O�O�O�O �O�O�O_ _=_$_6_ s_Z_�_~_�_�_�_�_ HO�_'o�_Ko2ooo�o ho�o�o�o�o�o�o�o #5Y@}dv �
o�����1� �*�g�N���r����� ���̏	���?�&� c�u����P���ϟ�� �ڟ�)��M�4�q� X�j�����˯���� �%�|��[���f� ������ٿ������� 3��W�i�Pύ�tϱ�p�Ϫ���7�d ���	���	�B�-�f�Qߌ�ߙ�%��߾�>�����у������� ����9�'�]�k�� ����S��������� ���;�}�b���+��� ������������C�i� :y�m[�� �� ?�3� CiW�{��� �/�///?/e/ S/�/��/�y/�/�/ ?�/+??;?a?�/�? �/Q?�?�?�?�?O�? 'Oi?NO`OO9OO�O �O�O�O�O�OAO&_eO �OY_G_i_k_}_�_�_ �__�_=_�_1ooUo Coeogoyo�o�_�oo �o	�o-Q?a �o�o��o���� �)��M��t��=� ��9���ݏˏ��%� g�L�����m����� ��ٟǟ��?�$�c�� W�E�{�i�������կ ���;�ů/��S�A� w�e���ݯ¿Կ���� ����+��O�=�sϵ� ��ٿc��ϻ������� '��Kߍ�r߱�;ߥ� ���߷�������#�e� J���}�k����� ����+�Q�"�a���U� C�y�g���������� '�����+Q?u c��������� 'M;q�� �a����// #/I/�p/�9/�/�/ �/�/�/�/?Q/6?H? �/!?�/i?�?�?�?�? �?)?OM?�?AO/OQO SOeO�O�O�OO�O%O �O__=_+_M_O_a_ �_�O�_�O�_�_�_o o9o'oIo�_�_�o�_ oo�o�o�o�o�o5 wo\�o%�!�� ����O4�s� g�U���y�������� '��K�Տ?�-�c�Q� ��u��������#��� ��;�)�_�M���ş ����s���o�ݯ�� 7�%�[�������K��� ��ſǿٿ���3�u� Zϙ�#ύ�{ϱϟ��� �����M�2�q���e� S߉�w߭ߛ߽��9� 
�I���=�+�a�O�� s����������� �9�'�]�K������ ��q���������5 #Y�����I�� ����1sX �!�y���� �9/0/�	/�Q/ �/u/�/�/�//�/5/ �/)??9?;?M?�?q? �?�/�??�?O�?%O O5O7OIOO�?�O�? oO�O�O�O�O!__1_ �O�O~_�OW_�_�_�_ �_�_�_o__Do�_o wo	o�o�o�o�o�o�o 7o[o�oO=sa �����3� '��K�9�o�]���� �̏������#�� G�5�k�������[�}� W�ş�����C��� j���3����������� ����]�B����u� c������������5� �Y��M�;�q�_ϕ� �ϥ���!���1���%� �I�7�m�[ߑ��ϸ� �ρ���}���!��E� 3�i�ߐ���Y���� ��������A���h� ��1������������� ��[�@�	sa �����! ���9o]�� ����/�!/ #/5/k/Y/�/��/� /�/�/?�/??1? g?�/�?�/W?�?�?�? �?	O�?Oo?�?fO�? ?O�O�O�O�O�O�O_ GO,_kO�O__�Oo_�_ �_�_�_�__oC_�_ 7o%o[oIoko�oo�o �_�oo�o�o3! WEg��o��o} ����/��S�� z���C�e�?����я ���+�m�R������ s�������ߟ͟�E� *�i��]�K���o��� ����ۯ��A�˯5� #�Y�G�}�k����	� ڿ������1��U� C�yϻ���߿i���e� ��	���-��Qߓ�x� ��A߫ߙ��߽���� ��)�k�P����q� ���������C�(� g���[�I��m����� ��	��� ������! WE{i���� ���	SA w���g��� �///O/�v/� ?/�/�/�/�/�/�/? W/}/N?�/'?�?o?�? �?�?�?�?/?OS?�? GO�?WO}OkO�O�O�O O�O+O�O__C_1_ S_y_g_�_�O�__�_ �_�_o	o?o-oOouo �_�o�_eo�o�o�o�o ;}obt+M '������U :�y�m�[�}���� Ǐ���-��Q�ۏE� 3�i�W�y�{���ß� �)�����A�/�e� S�u�˟�¯����� ���=�+�a����� ǯQ���M�˿�߿� �9�{�`ϟ�)ϓρ� �ϥ��������S�8� w��k�Yߏ�}߳ߡ� ����+��O���C�1� g�U��y�������� �����	�?�-�c�Q������������$S�ERV_MAILW  ��������OUTPUT�����@��RoV 2w�  ��� (��I��S�AVE��TOP�10 2#	 d ����� �'9K]o �������� /#/5/G/Y/k/}/�/ �/�/�/�/�/�/?? 1?C?U?g?y?�?�?w��{YPf��FZN_CFG w���W�1?GRP 2�7t� ,B   A�'@��D;� B�(@�  B4��RB21VHELL�2	w�r6 �7�7�O�K%RSR�O�O�O�O�O_ �O3__W_B_T_�_x_��_�_�_�_�_on�  ��RoKoX]o+bio ��eoL�b�`�bg3b2���dultm�bRFHK ;1
`K �o 0YTfx� �������1��,�>�P�LLOMM �`O��QBFTOV_ENB��+r��bOW_REG_�UI����IMIO/FWDL����*E^��WAIT���i��2����*�T�IM���T�V�A��+���_UNI�T����r	LCڀT�RY�r��M�ON_ALIAS� ?e��2 he ���!�3�E�S���v� ������W�Я���� �ï<�N�`�r���/� ����̿޿𿛿�&� 8�J���[πϒϤ϶� a��������"���F� X�j�|ߎ�9߲����� ���ߥ��0�B�T��� x������k����� ��,���P�b�t��� ��C����������� (:L^	��� ��u� $6 �Zl~��M� ���� /2/D/V/ h//�/�/�/�/�// �/
??.?@?�/d?v? �?�?E?�?�?�?�?O �?*O<ONO`OrOO�O �O�O�O�O�O__&_ 8_J_�On_�_�_�_O_ �_�_�_�_o�_4oFo Xojo|o'o�o�o�o�o �o�o0B�oS x���Y��� ���>�P�b�t��� 1�����Ώ��򏝏� (�:�L���p������� ��c�ܟ� ��$�Γ��$SMON_D�EFPROG �&���N�� &*SY�STEM*+�o�����?=�RECALL ?}N�� ( �}
x�yzrate 1�1 =>169.�254.��120:19636 ��`ĥ�����}!��24��ǯٯj�|����!�:copy f�rs:order�fil.dat �virt:\tm?pback\5�`�����}1��mdb:*.*��ѿJ�`ݿnπϒ�%�5x��:\3ϴ�E�G�`���,��}6��a���� B���r߄�ߩ���D� _�����'���K��� n����8�E����� ���#ߴ���Y�j�|� ���߳�<������� �1���U�fx��� ��B������-� �Q��t����5 GY��/!�3�E� 7/�o/�/�/�5/G/ Y/�/�/?!/3/�/�/ h?z?�?�/�/C?U?�? �?
O?/?�?�?dOvO �O�?�??OQOcO�O_ O+O�O:_�Or_�__ �O;_�___�_oo'_ �_�_�_no�o�o�_Lo Io[o�o�o#o�o�o �oj|��o�oEW ���1��f� x�����A�S���� ��-���я�t��� ����=���a����� )���8�ߟp������� N�K�]�� ��%�̯ ɯۯl�~�������> ������!�οW h�zόϟ����� ��
�/��S�d�v� �ߛ���6�M�c���� �+���O���r�����$SNPX_A�SG 2������� 7 0��%������  ?���PAR�AM ��^�� �	��P�������1������OFT_KB_CFG  ������OPIN_S_IM  ��,�����������RV�NORDY_DO�  6�b���QSTP_DSBv��,���SR }�� � &0��Q����G�TOP_ON_ERR�����|PTN z��� �A��RING_PRM����VCNT_G�P 2x�.���x 	
	���0�T��VD� RP 1�/�E��7 �������/ /1/C/U/g/y/�/�/ �/�/�/�/�/	??-? ??Q?c?�?�?�?�?�? �?�?�?OO)OPOMO _OqO�O�O�O�O�O�O �O__%_7_I_[_m_ _�_�_�_�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /Ahew��� �����.�+�=� O�a�s���������͏ ����'�9�K�]� o���������ɟ۟� ���#�5�G�Y���}� ������ůׯ���� �F�C�U�g�y����� ����ӿ��	��-��?�Q�c�mPRG_�COUNTW�眯��ENB���M���Y���_UPD �14T  
 xϣ���/�X�S�e� wߠߛ߭߿������� �0�+�=�O�x�s�� ������������ '�P�K�]�o������� ����������(#5 Gpk}���� � �HCU g������� � //-/?/h/c/u/ �/�/�/�/�/�/�/? ?@?;?M?_?�?�?�? �?�?�?�?�?OO%O 7O`O[OmOO�O�O�O���_INFO 1=����P	 �O__@_+Y�@l�@I�l�?Z�F_-S��̵��5A�u�9	�]�ƿ��@�K]A����@CP A?!" ?�nn_�A� D5Oy����C����($6�T5�+���Q� �8�h�Ca����.~:��1�５���YSDOEBUG������@�d��
`SP_PA�SS��B?kL_OG �Fї  �@�X�O � ����AUD�1:\Hd�NIb_M�PCNm���o�o���a�o ���fSAV Qi��2Qqa�b��E�hSV�kT�EM_TIME �1Qg� 0
�������Z���^s�MEMBK  ����q`qo�� ��X|��� @ ��C�"�G�W��dz�����a 2[@}q��я���/s���1�C�U�g�y� � {�����ß՟�����/�i�e>�c�u��� ������ϯ���� )�;�M�_�q���������\uSK�p�x���������1�@|���2,�W�AW΀A Tý�i��Ϧ�(��#!������� ���<�-�  �-���0��s߅ߗߋ�X����������(��@$,�P�D�t���� ����������(�:� L�^�p��������������T1SVGUNwSPD2e 'e����2MODE_LIM �vvq b2��2��Qm���ASK_OPTI�ON`�y aS_�DI+`ENB  �b�esBC2_?GRP 2ܵc|r�[R��C������BCCFG ��7| (��`M_VAf� w������/ //R/=/v/a/�/�/ �/�/�/�/�/??<? '?`?K?�?�?8Ձ<�? �?�?�?p?�?+OOOO :OsO~�O�th@�O�O �O�O�O	_�O-__=_ ?_Q_�_u_�_�_�_�_ �_�_o)ooMo;oqo _o�o�o�o�o�o�o�h �03EW�o{ i������� ��A�/�e�S�u�w� �������я���+� �;�a�O���s����� ͟��ݟߟ�'��K� c�u�������5�ۯ ɯ����5�G�Y�'� }�k�����ſ��տ׿ ���C�1�g�Uϋ� yϛ��ϯ�����	��� -��=�?�Q߇�u߫� a����������;� )�K�q�_����� �������%��5�7� I��m����������� ����!E3iW �{����� ��#5Sew�� �����//� =/+/a/O/�/s/�/�/ �/�/�/?�/'??K? 9?[?�?o?�?�?�?�? �?�?�?�?OGO5OkO !�O�O�O�O�OUO�O �O_1__U_g_y_G_ �_�_�_�_�_�_�_�_ 	o?o-ocoQo�ouo�o �o�o�o�o�o) M;]_q��� �O���%�7��[� I�k������Ǐُ�� ���!��E�3�U�W� i�����ß���՟� ���A�/�e�S���w� ��������ѯ���+� �C�U�s�����������˿�߿���3���$TBCSG_G�RP 2���  �3�� 
 ?�   ^�p�Zϔ�~ϸϢϴ�@�����$�7�>�E̿d0 �S�?�3�	 HCA��"�>l�"�CS�BpVߙ�c�u߇����B�$�>������"�Bl����)�A������G�"�;�B�)�+�Q�G��$_��A3�"�Q���T��Ѩ��@����� '�:���e���M�_�x������?�ff��� ��	V3.0}0V�	mt2 * 2�$��<23�G�� [ -\  q��7�+J2>�E����CFG !��eO� R��
����0� 0Vd�d�u� �����/// P/;/t/_/�/�/�/�/ �/�/�/??:?%?^? I?�?m??�?�?�?�?  OOV�p�O/OAO�? tO_O�O�O�O�O�O�O �O_(_:_L__p_[_ �__�_�_3���_�� �_ooIo7omo[o�o o�o�o�o�o�o�o 3!WEgi{� �������-� S�A�w�e�����m�ŏ ׏������=�+�a� O���s�����͟ߟ�� ���9�'�]�o��� ��M�����ۯɯ�� ��5�#�Y�G�}�k��� ����׿ſ����� C�1�S�U�gϝϋ��� ������	����?�� W�i�{�%߫ߙ߻߽� �����)��M�_�q� ��A��������� �%���5�[�I��m� ��������������! E3iW�{� �����/ ?AS�w��� ����/��O/=/ s/a/�/�/�/�/�/�/ ??�/%?K?9?o?]? �?�?�?�?�?�?�?O �?!OGO5OkOYO�O}O �O�O�O�O�O_�O1_ _U_C_y_g_�_�_�_ �_�_�_�_o	o+o-o ?ouo��o�o�o[o�o �o�o;)_M ����w��� ��7�I�[��'��� �����ُǏ���� 3�!�W�E�{�i����� ����ß�����A� /�e�S�u��������� �ѯ���o1�C��o ����s�����Ϳ��ݿ ��'�9�K�	�ρ� oϥϓ��������Ϲ� #��3�5�G�}�kߡ� ���߳��������� C�1�g�U��y��� ������	���-��Q� ?�a���u���%�W��� ������M;q _������� #%7m� �]����/� /!/3/i/W/�/{/�/ �/�/�/�/?�//?? S?A?w?e?�?�?�?�? �?�?�?OO=OOO�� gOyO�O5O�O�O�O�O �O�O_9_'_]_o_�_ �_Q_�_�_�_�_�_�^�  %`)c �)f=o)b�$TBJ�OP_GRP 2�"�U� _ ?�)f	Ub�\c$cl��P��pJ�`��xe  � �� � ��`�)d� @%`tb	 ��CA��f��S�C��_)eta�b3�33�f�oz=�_��CS�?��Y�1ru`B�;pp�gLWw�o�o?�a�u�ޜz<؄-r��a��u=�)eB��w?C�  D�a�o�#�-�;��B9l�`2u�ff�n�&)eAЇ��w���>��ͭ�����;�ǎ���@fff���b�]���A���������9�ˌ�X��@�o�폎������%��ɟۛ;������@�o��� {����9�1�g�Y�C� Q������E�ϯ�ӯ ��@��կ_�y�c�Pq���пct�)f���	V3.00�zcmt2��*��yd$a)�4� �F� G9| �G�v�G�/��G�� H�@�H,�H.���HC� HYA@�Hn��H�� �H�� H�Y@�H�`H����H�c�H��H̿�H�nD��G G.A �GKm Gh� �G��G�x��G��G����G�:�G�Ѐ�G�f�G����G��\��H
�_�H��H���H @�H'��d�ր=L��=#�
������)bQ3o�+�)f/��?�߀f�d�RcESTPARS�hn`�RcHR��ABLEW 1%ci�)d�_�D� �@$�_�B_�_�(g0a_�	_�E
_�_ؾ�)a_��_�_�����RD	I��ma�����������O������������S��kc  I���������� *<N`r��� ����Hm���� lb��C,�>�P�b�� �2�D�V�h��)N�UM  �U*ma�`1` ������_CFG &�+��a@U`IMEBF_TT�Ѻkc��T&VER�Uj&�T#R 1'��' 8&�)b$`�! �PN  �/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? <OO)OrOMO_OuO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_4oo!ojo EoWomo{o�o�o�o�o�җ!_!�&@�%���MI_CHAN�`' �% .sDBGLVL`'�%��1p�ETHERAD �?���p�/���o�o��y�1pRO�UT~ !�!��t��|SNMAS�Kyx�#�q255.?��=�O�a�Á��OOLOFS_D�I���ecyORQCTRL (�+��0�ߍTΏ��'� 9�K�]�o��������� ɟ۟����#�3�͏�V�E�z�~�PE_D�ETAIWx��PG�L_CONFIG� .)"!���/cell/$C�ID$/grp1�~�����*�<��� �g�y���������P� ���	��-�?�οc� uχϙϫϽ�L�^��� ��)�;�M���q߃� �ߧ߹���Z����� %�7�I��������������M}n��!� 3�E�W�i��k���p��m���������  g�DVhz��- ����
.� Rdv���;� ��//*/�N/`/ r/�/�/�/�/I/�/�/ ??&?8?�/\?n?�? �?�?�?E?�?�?�?O "O4OFO�?jO|O�O�O �O�OSO�O�O__0_ B_�Of_x_�_�_�_�_��_͠�User View ��}}1234567890oo'o9o�Ko]oed�`£�o���Y2�Yb_�o�o�o�o !�o�o�R3�oo �����(��n4^#�5�G�Y�k�}�����n5�׏���@��1���R��n6Ə ��������ӟ�D���n7z�?�Q�c�u����������n8.�����)�;�M���n�t� �lCamera�Z꯳�ſ׿������E��7�I� [�ouχϙϫϽ���ŉ  ���i���1� C�U�g�y� ϝ߯��� �����	��-�?�f����]y�ߋ����� �����	��-�x�Q� c�u�������R�d�� B���	-?Q�� u�������� ��d��˰ew ����f��/ R+/=/O/a/s/�/, ��y�/�/�/�/?? )?�M?_?q?�/�?�? �?�?�?�?�/d�-��? ;OMO_OqO�O�O<?�O �O�O(O__%_7_I_ [_Od���O�_�_�_ �_�_o�O%o7oIo�_ moo�o�o�o�on_�W9So,>Pb 	os��Qo������(�:�ɪ	��0 �u���������Ϗv ����;�M�_�q� ����<�N�����9��  ��$�6�H��l�~� ��۟��Ưد���� ����ۥ�Z�l�~��� ����[�ؿ���G� � 2�D�V�h�z�!�[�n� ���������� �ǿ D�V�h߳όߞ߰��� ���ߍϟ���}�2�D� V�h�z��3߰����� ���
��.�@�R��� ��F����������� ����.@��dv ����e��Ų+U 
.@Rd� ������//<*/�  �	Y/ k/}/�/�/�/�/�/�/x�/?;   // 7/U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o�#<  
� (  ��M ( 	  �o�o�o�o�oC 1SUg����t��j?: �y *�<�N��r������� ��̏������a� >�P�b�t�����ߏ�� Ο��'���(�:�L� ^����������ʯܯ � ��$�k�}�Z�l� ~�ů����ƿؿ��� C� �2�Dϋ�h�zό� �ϰ���	�����
�Q� .�@�R�d�v߈����� ������)���*�<� N�`�߄������� ������&�m�J�\� n�������������� 3�E�"4F��j| ������ S0BTfx�� ����//,/ >/P/���/�/�/� �/�/�/??(?o/L? ^?p?�/�?�?�?�?�? �?5?O$O6O}?ZOlO�~O�O�O�O�?�p@ A�B�O�O_�C�G��`��#frh:�\tpgl\ro�bots\m10�iaAS_8l.xml�Oe_w_�_�_�_��_�_�_�_on�� o>oPoboto�o�o�o �o�o�o�oo: L^p����� �� ��6�H�Z� l�~�������Ə؏� ����2�D�V�h�z� ������ԟ���� 	�.�@�R�d�v����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶���������� XVA |�O+P<< )P ?���A���9�[� ��oߑ߿ߥ������� ���=�#�E�s�Y������������6��$TPGL_OUTPUT 1	A�	A !� -�B�T�f�x������� ��������,> Pbt�������-�!Є��2345678901 );M_g�2 ��������@/0/B/T/f/�}p/ �/�/�/�/�/x/�/? (?:?L?^?p??~?�? �?�?�?�?�?�?$O6O HOZOlOOO�O�O�O �O�O�O�O
_2_D_V_ h_z__�_�_�_�_�_ �_�_�_.o@oRodovo �o o�o�o�o�o�o �o<N`r� .������� "�J�\�n�����*����ȏڏ�������} �F�X�j�|��������@#�՟�)� ( 	 ��
�@� .�d�R���v������� �Я���*��N�<� ^���r�����̿��� ޿ ���J�8�n����8�vϨϺ͒��� �����$��
��U�g� �sߝ�w߉�����C� �����Q�c�=�� ���߁���i���� ��;�M���5�����/� ��������_�q�7 I��QYk�� %����3 i{���K�� ��///�/e/w/ /�/�/�/�/�/A/�/ ?+?�/O?a?;?M?�? �/?�?�?y?�?O�? OKO]O�?aO�O-OO �O�O�O�O_oO�OG_ �O3_}_�_i_�_�_#_ �_�_o�_1oCooOo yo�_�_�o�o[o�o�o �o�o-?�ocu�a�������)�WGL1.XM�L��(��$TPOFF_LIM ��|�����6��N_SV>�  ���P�P_MON7 2��R������22�STRT?CHK 3��P��C�9�VTCOM�PATe��T�VW�VAR 4��\�i� Ə *��I���:�_DE�FPROG %���%MAINo  TLd�T1A��3�_DISPLA�YE���Z�INST�_MSK  ��� ��INUSE9R叜�LCK�QUICKME{���Z�SCRE1������tps�c���L�Q�P�b�_�f�ST�P�RAC�E_CFG 5����I�	3�
�?���HNL 2!6i�b�ѡ� ?�� �)�;�M�_�q��������ITEM 27�� �%$12�34567890<ؿ�  =<��<�"�  !(�0�<��u�3�ֿ���� ����0���T�f�/ߊ� J߮�Z߀������ 4�>߸�b��4�F�� j�������l������ ��^������*�x� ��������6�H� l�,��Pb��x�� <� �D�( �4���N�� ��@ /dv�/ $/�~/�/��//*/ �/N/?r/2?D?�/Z? �/�/�??�?&?�?�? ~?n?�?�?�?�?0O�? �O�O�O"O�OFOXOjO �O�O:_`_r_�O~_�O __�_�_T_o&o�_ 2o�_�_�o�_�oo�o �o>o�obo�o=�oX �oh���(: L�p�B�T��x� �� �����6���� l������k�Ə��� ���� �ҟD�V�����S��8��$�� 3 ��$� ɡ{�r�
 ������ү~S�UD1:\߬���6�R_GRP� 19Ż� 	 @{�*�<�&�@\�J���n�������� ˿ٺ��߯��'��?�  B�T�>�t� bϘφϼϪ������� ��:�(�^�L߂�p��߸�	�����4��SCB 2:@� -�*�<�N�`�r�������*�UTORIAL ;@��Ư�/�V_CON?FIG <@�ġ�x�¯d��OUTP�UT =@�U���p��������� �� 2DVhz �R�������  2DVhz� ������
// ./@/R/d/v/�/��/ �/�/�/�/??*?<? N?`?r?�?�?�/�?�? �?�?OO&O8OJO\O nO�O�O�?�O�O�O�O �O_"_4_F_X_j_|_ �_�O�_�_�_�_�_o o0oBoTofoxo�o�o �_�o�o�o�o, >Pbt���o� �����(�:�L� ^�p��������ʏ܏ � ��$�6�H�Z�l� ~�����>�P������ ��(�:�L�^�p��� ��������ܯ� �� $�6�H�Z�l�~����� ��ůؿ���� �2� D�V�h�zόϞϰ��� ӿ����
��.�@�R� d�v߈ߚ߬߾����� ����*�<�N�`�r� ������������ �&�8�J�\�n����� ������������" 4FXj|��� �����0B Tfx����� ��//,/>/P/b/ t/�/�/�/�/�/��/ ??(?:?L?^?p?�?��?�?�?�?������?�?�1�?&Oɟ JO\OnO�O�O�O�O�O �O�O�O_"_�/F_X_ j_|_�_�_�_�_�_�_ �_oo0oA_Tofoxo �o�o�o�o�o�o�o ,=oPbt�� �������(� 9L�^�p��������� ʏ܏� ��$�6�G� Z�l�~�������Ɵ؟ ���� �2�C�V�h� z�������¯ԯ��� 
��.�?�R�d�v��� ������п����� *�<�M�`�rτϖϨ� ����������&�8� I�\�n߀ߒߤ߶��߀�������"�4�C���$TX_SCRE�EN 1>�5w�0�}�C�@���������u� 2Ft�!�3�E�W�i�{� ������������� ��/��Sew�� �$�H�+ =O������ ��V/z'/9/K/ ]/o/�/��//�/�/ �/�/?#?�/�/Y?k? }?�?�?�?*?�?N?�?�OO1OCOUO�?yO��$UALRM_M_SG ?c��p� qOFګO�O�O�O __6_)_;_Y___�_��_�_�_�_�ESEV7  �M
f�BECFG @c�m�  F�@�  A:a   ;B�F�
 �_M� c�moo�o�o�o�o�o��o�o!/waGR�P 2A k 0�F�	 Woy�@I�_BBL_NOT�E B jT��lM�h�O��,`�rDEFPR�O�@%�K (%�MAINz�}% �_��?�*�c�N��� r��������̏��{�FKEYDATA� 1Cc�cpp 	/gF�fi�{�R�������,(���F��(POINT �ER��  OO�K O�C�ҐND�IRECTD�F� CHOICE]p���TOUCHUP����ȯ�ӯ��� 4�F�-�j�Q��������Ŀ������ω����/frh/g�ui/white�home.png�)�g�yϋϝϯπ>@�pointR���`����+ߺ�  A�look����k�}���ߡ߳�B�indirec�������#�|5�@�choicQ�@o������@�touchup_�@����+�=���@�arwrg��w��� ������F�����  $6H��l~�� ��U�� 2 D�hz���� �c�
//./@/R/ �v/�/�/�/�/�/_/ �/??*?<?N?`?7� e?�?�?�?�?�?�?�/ 
OO.O@OROdO�?�O �O�O�O�O�OqO�O_ *_<_N_`_r__�_�_ �_�_�_�__o&o8o Jo\ono�_�o�o�o�o �o�o�o�o"4FX j|����� ���0�B�T�f�x� �������ҏ���� ��,�>�P�b�t���� ����Ο��������:�L�^�p�����/�����:����ʯܯ�Ư�"���,�S��w�^����� ��ѿ������+�� O�a�Hυ�lϩϻϢ� �������'�9� �]� D߁ߓ�r?�������� ��� �5�G�Y�k�}� ���0���������� ���C�U�g�y����� ,���������	- ��Qcu���: ���)�M _q����H� �//%/7/�[/m/ /�/�/�/D/�/�/�/ ?!?3?E?�/i?{?�? �?�?�?R?�?�?OO /OAO�?eOwO�O�O�O �O�O���O__+_=_ O_VOs_�_�_�_�_�_ �_n_oo'o9oKo]o �_�o�o�o�o�o�ojo �o#5GYk�o ������x� �1�C�U�g������ ����ӏ������-� ?�Q�c�u�������� ϟ�󟂟�)�;�M� _�q��������˯ݯ ����%�7�I�[�m� ������ǿٿ������@���@���:�L�^�6��ϒ�l�,~���v��� �����A�(�e�w� ^ߛ߂߿��߸����� �+��O�6�s�Z�� ����������O'� 9�K�]�o��������� ����������5G Yk}���� ���1CUg y��,���� 	//�?/Q/c/u/�/ �/(/�/�/�/�/?? )?�/M?_?q?�?�?�? 6?�?�?�?OO%O�? IO[OmOO�O�O�ODO �O�O�O_!_3_�OW_ i_{_�_�_�_@_�_�_ �_oo/oAo�eowo �o�o�o�o�_�o�o +=O�os�� ���\���'� 9�K��o��������� ɏۏj����#�5�G� Y��}�������şן f�����1�C�U�g� ����������ӯ�t� 	��-�?�Q�c�򯇿 ������Ͽ�󿂿� )�;�M�_�q� ϕϧ� ��������~��%�7ߠI�[�m��V`��}�V`�����@���ݦ������,�� 3���W�>�{��t�� �����������/�A� (�e�L����������� ���� =$a sRo������  �'9K]o� ������� #/5/G/Y/k/}//�/ �/�/�/�/�/?�/1? C?U?g?y?�??�?�? �?�?�?	O�?-O?OQO cOuO�O�O(O�O�O�O �O__�O;_M___q_ �_�_$_�_�_�_�_o o%o�_Io[omoo�o �o2o�o�o�o�o! �oEWi{��� ������/�6 S�e�w���������N� �����+�=�̏a� s���������J�ߟ� ��'�9�K�ڟo��� ������ɯX����� #�5�G�֯k�}����� ��ſ׿f�����1� C�U��yϋϝϯ��� ��b���	��-�?�Q� c��χߙ߽߫����� p���)�;�M�_��� ������������p�����p����,�>��`�r�L�,^��V������ ����!EW>{ b������ �/S:w�p �����//+/ =/O/a/p�/�/�/�/ �/�/�/�/?'?9?K? ]?o?�/�?�?�?�?�? �?|?O#O5OGOYOkO }OO�O�O�O�O�O�O �O_1_C_U_g_y__ �_�_�_�_�_�_	o�_ -o?oQocouo�oo�o �o�o�o�o�o); M_q��$�� �����7�I�[� m���� ���Ǐُ� ���!��E�W�i�{� ������ß՟���� �/���S�e�w����� ��<�ѯ�����+� ��O�a�s��������� J�߿���'�9�ȿ ]�oρϓϥϷ�F��� �����#�5�G���k� }ߏߡ߳���T����� ��1�C���g�y�� �������b���	�� -�?�Q���u������� ����^���);hM_6�a�6�����������,�� 7[mT�x� ����/!//E/ ,/i/{/b/�/�/�/�/ �/�/�/??A?S?2� w?�?�?�?�?�?���? OO+O=OOOaO�?�O �O�O�O�O�OnO__ '_9_K_]_�O�_�_�_ �_�_�_�_|_o#o5o GoYoko�_�o�o�o�o �o�oxo1CU gy����� ���-�?�Q�c�u� �������Ϗ��� ��)�;�M�_�q���� ����˟ݟ����%� 7�I�[�m����h?�� ǯٯ�����3�E� W�i�{�����.�ÿտ ����Ϭ�A�S�e� wωϛ�*Ͽ������� ��+ߺ�O�a�s߅� �ߩ�8��������� '��K�]�o���� ��F��������#�5� ��Y�k�}�������B� ������1C�� gy����P� �	-?�cu@�����������������/-�@/R/,&, >?�/6?�/�/�/�/�/ ?�/%?7??[?B?? �?x?�?�?�?�?�?O �?3OOWOiOPO�OtO �O�O���O�O__/_ A_Pe_w_�_�_�_�_ �_`_�_oo+o=oOo �_so�o�o�o�o�o\o �o'9K]�o ������j� �#�5�G�Y��}��� ����ŏ׏�x��� 1�C�U�g��������� ��ӟ�t�	��-�?� Q�c�u��������ϯ �󯂯�)�;�M�_� q� �������˿ݿ� ��O%�7�I�[�m�� ���ϵ���������� ��3�E�W�i�{ߍ�� ������������/� A�S�e�w���*�� ����������=�O� a�s�����&������� ��'��K]o ���4���� #�GYk}� ��B���// 1/�U/g/y/�/�/�/ >/�/�/�/	??-???��A;�����j?|?�=f?�?�?�6,�O�?�OO�? ;OMO4OqOXO�O�O�O �O�O�O_�O%__I_ [_B__f_�_�_�_�_ �_�_�_!o3o�Woio {o�o�o�o�/�o�o�o /A�oew� ���N���� +�=��a�s������� ��͏\����'�9� K�ڏo���������ɟ X�����#�5�G�Y� �}�������ůׯf� ����1�C�U��y� ��������ӿ�t�	� �-�?�Q�c��ϙ� �Ͻ�����p���)� ;�M�_�q�Ho�ߧ߹� ���������%�7�I� [�m��������� �����!�3�E�W�i� {�
������������� ��/ASew� ������ +=Oas��& ����//�9/ K/]/o/�/�/"/�/�/ �/�/�/?#?�/G?Y? k?}?�?�?0?�?�?�? �?OO�?COUOgOyOЋO�O�O���K�>������O�O �M�O _2_V,oc_ o�_n_�_�_�_�_�_ oo�_;o"o_oqoXo �o|o�o�o�o�o�o �o7I0mT�� �������!�0O E�W�i�{�������@� Տ�����/���S� e�w�������<�џ� ����+�=�̟a�s� ��������J�߯�� �'�9�ȯ]�o����� ����ɿX�����#� 5�G�ֿk�}Ϗϡϳ� ��T�������1�C� U���yߋߝ߯����� b���	��-�?�Q��� u��������� ��)�;�M�_�f�� ������������~� %7I[m���� ����z!3 EWi{
��� ����///A/S/ e/w//�/�/�/�/�/ �/?�/+?=?O?a?s? �??�?�?�?�?�?O �?'O9OKO]OoO�O�O "O�O�O�O�O�O_�O 5_G_Y_k_}_�__�_��_�_�_�_oo�$�UI_INUSE�R  ����@a� �  o$o_MENHIST 1D@e�  �( M`��(/�SOFTPART�/GENLINK�?current�=menupage,153,1_o0�o�o�o�'�o�n71�oSew��Qy)�eedit�bMAINB���p��,�`422��]�o�����4�e,�2�oޏ�����R� �>�P�b�t�����'� ��Ο�������:�@L�^�p��������4� �a4�ѯ�����+� .�O�a�s�������8� Ϳ߿���'϶�ȿ ]�oρϓϥϷ�F��� �����#�5���Y�k� }ߏߡ߳�B�T����� ��1�C���g�y�� ����אָ����	�� -�?�Q�T�u������� ����^���); M_������� �l%7I[ ������� z/!/3/E/W/i/� �/�/�/�/�/�/���� ?/?A?S?e?w?z/�? �?�?�?�?�?�?O+O =OOOaOsO�OO�O�O �O�O�O_�O'_9_K_ ]_o_�__�_�_�_�_ �_�_o�_5oGoYoko }o�oo�o�o�o�o�o �/
?CUgy� ��o����	�� ��Q�c�u������� :�Ϗ����)��� M�_�q�������6�H� ݟ���%�7�Ɵ[� m��������D�ٯ�����!�3���$�UI_PANED�ATA 1F����i� � 	�}  f�rh/cgtp/�flexdev.�stm?_wid�th=0&_height=10�����ice=TP&�_lines=3���columns�=4��fon��4�&_page=d�oub��1E�!v)�  rim��  z�(�:�L�^�pς� 鿔ϸϟ����� �� ��6��Z�l�Sߐ�w����߭���!v� ��    � �v"�FR�H/VISION�/VRFRMN.STM?_imӰ�only=1ǰi�ltershow�n��A�ed=1 亿̿2���ual ���$��������� /���S�:�w���p��� ����������+ OaH����k� �����%x I��m���� .���!//E/W/ >/{/b/�/�/�/�/�/ �/�/?/?��e?w? �?�?�?�??�?VO O+O=OOOaOsO�?�O ~O�O�O�O�O�O_�O 9_K_2_o_V_�_�_�_ �_<?N?�_o#o5oGo Yo�_}o�oO�o�o�o �o�oto1Ug N�r����� 	���?�&�c��_�_ �o����Ϗ���X� )��oM�_�q������� �˟ݟğ��%�7� �[�B��f������� ٯ���������E�W� i�{������ÿ6�� ����/�A�SϺ�w� ^ϛςϿ��ϸ����� �+��O�6�s߅�l� ���.�������'� 9��]�o�⿓��� ������T����5�G� .�k�R����������� ������C����}�T������){��8J \n������ ��/�4//X/j/ Q/�/u/�/�/�/�/x�������$UI_P�OSTYPE  ���� �	 �/K?2QU�ICKMEN  �);8?N?0RE�STORE 1G���  '��/���?�3�?��m�?O+O=OOO aOO�O�O�O�O�OpO �O__'_9_�?F_X_ j_�O�_�_�_�_�_�_ o#o5oGoYokoo�o �o�o�o�o�_�o�o zoCUgy�.� ������-�?� Q�c��������� ����)�̏M�_� q�����8���˟ݟ� ���� �2���m�� ������X�ٯ���� !�3�֯W�i�{������Y7SCREi0?�n=u1sc��0u2ڴ3ڴ4�ڴ5ڴ6ڴ7ڴ8�ڱ��TAT%=� �}3��:USER�����Ӵksܳm�3�m�4m�5m�6m�7�m�8m�0NDO_?CFG H);d �c0PD�W��None\2�N�_INFO 1�I���{00% ���x�
�K�.�o߁� dߥ߷ߚ��߾������5�G�*�k�R<��O�FFSET L)9�x�@��0H��� ��������(�U�L� ^���b����������� ��$6��~?��p�
����UFRAME  @������RTOL_�ABRT���E�NB GRP �1M�9z1Cz  A�ec��cu ������h0�U/��MSK � 2�N��%���%Rs/ _'EVN2$�ƈ&v��2N��
 h���UEV!�td:\event_user\w/F� C7�/�B�F<��!SP�!�'sp�otweld=!C6????�0b$!b/�/�?�?�7!�? �?�?OAO�?�?wO"O �OFOXOjO�O�O_�O �O�OO_>_s__0_f_ �_�_�_�_�_o�_9o Ko�_o�o,o�oPobj~�&WRK 2OX�F�8�o	 �o @R-v�c�� �����*��N� `�;�����q���̏���ݏ���$VARS_CONFI���P�� FP@����CCRG��SP��Z@�9�D��B�BH�p����Ce���їϑ?�ᐶU�MRK2Y��)B�	��C�X��1: SC13?0EF2 *3�7��@����ch �5�B����A@��C�Ȑ� ��� ��9���ȯ�����"���ӑ��	�Z���� B��� u���z����᯾��� �Ϳ��*��'�`� ��Aϖρϓ������\�X�TCCc�ZR��4��pa��'�G�F,��![�� ��a 2345678901q�y�'9�n���n߰ߘ#����j�$����B��Ӗ ��ϑ?:�o=L{�� !p� �p��ia/[�� �Ԇ���������� )�;�(�:�q��p��� ���������%� I�[�H���{���������"�S�SELE�C�$!?�AVIoA_WO�`\T)�_ff,		��= �;G�P ��R'	�RTSYN'CSE�j��n�e�WINURL ?u��R����� //"�ISI�ONTMOU�/ ��*%c�]S۳��S۵@/� �FR:\,#\D�ATAs?MЄ� wMCk&LOGx/   UD1k&�EX�/��' ?B@ ���"�!�DESKTOP�-MC6FJ6K��/�#?%?�le �� n6  �����f�"�� -��N5K�   =���w1��t0� }�(TRAIN�/hH҆2�bd�3pw5>{4 #`�"'(:��^]� (���9 M��OO+O=OOO�O sO�O�O�O�O�O�O�O�_$(STAT _'� �z�b_t_�_�hq$�_�_'%_GES#�`]���0 �
����R�WHOMI}NV aS۾�`��b"���C�ז�&�WJMPERR� 2b]�
   =�jho^l��o�o�o �o�o�o�o.<�m`r�S_� R�EV cO^#�LEXr�Td7��1-e�_�VMPHASE � j���&�O�FFo_ENB � \�	P2R$e/SۿN��c|3�@:�`Q�u����?s33�4�1K� g�']g�t�g��&�S`�hWm�3�\C*��J��������81��_�
�A/�4��/�7k� C9�qA�т�/�Q�� S�4�0�3��o�=�,������5ǟ[@3�B�7Ϋ�o����A�A�;2C%���c_������]�s�����^����9¸�+��3�����%����(��}��+}�eC�����A�W������ݔ�&��I�J.+c����v{)Kw@��#߯Կ�1������Y�*"H���P*�g���/�y���i��'�=σ�xϺ�%�B�L��s��#)���
���2�ÿ��������B�ՠ��7�4o��*	H�C���E���_�T�XB��krCI��a#��ܫC%r�ا������M�B�;C�6��E�����+�eB�5���)�����C߀8�X��߄�� [��������3� ���i�^�p������ ������� /�!S� Hw�����y��� ���+=2a��_q��ÅTD�_FILTES`i��[ Է��P�� <//'/9/K/]/o/ �/�/�/6��/�/�/ ??,?>?P?b?t?�Y�SHIFTMENoU 1jWm<�|%��?�t�?�?O�? �?EOO.O{OROdO�O �O�O�O�O�O�O/__�	LIVE/S�NAP#Svsf�liv�~A_�^�PION &�U^PdRmenuz___��_�_�r�5G�kΉ�ֈ9MOG�l�~�z�łZDdm��a<�ۀ �P�$WA�ITDINEND�  �U��#bxfO9K-��oOUT�o�h�S�o�iTIM�e���lGo}�o2{��oz�oz�o�hREcLE�.��hTM^{�d�xc_ACT�WP-���h_DATOA n΅�%�_xB��6�rRDIS^P~�~�$XVRa�o9n�$ZAB�C_GRP 1p.[k ,2J��=�Qa�pVSPT qq9m�À�
�Z��_��Z)�?�އD/CSCH`r#������IPbs[o�!۟���؊MPC�F_G 1t������0�� O����u췙��p��� �	?���o`�  �?Ӡ2?�k��1�?�ɾ�����4/6��u��D5Oy����C���?����<�� ��>%��6�����u=�������ί�> ����Ɇ�����˿� � �8�h�Ca����.~:��1�����۸� #�&� �2�H�Vπ��,�>��0V�h��� ��`v����_CYL�IND�w(� ��� ,(  *E�V��B��fߣ��� ��������?�  ��D�+�=�z�ߞ� ��������g����@�'���v����̞�29x �� �=��� ?��	��-=��`���zA��SPHERE 2y%����*���� X�kFX��| ����///e wT/�x/_/q/�/���/�/�/��ZZ�v �f