��  	c4�A��*SYST�EM*��V9.1�0214 8/�21/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP6fBI�IZ@!�LRM_RECO�"  � ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� ."��!_I�F� � 
$_ENABL@C#T� P dC#U5K�!CMA�B �"�
� �OG�f 0CUR�R_D1P $Q3LI�N@S1I4$C$AU�SOd�APPI�NFOEQ/ 9�L A ?1�5�/ H �7�9EQUIP �2�0NAM� ���2_OVR�?$VERSI� �����0COUPL}E,   $�!;PPV1CES C �G1�!�PR0�2�	 � $SO{FT�T_IDB�TOTAL_EQ2� Q1]@NO`BU �SPI_INDE�]uEXBSCRE�EN_�4BSI�G�0O%KW@P�K_FI0	�$THKY�GPA�NEhD � DU/MMY1d�D�!RU4 Q!RG1R��
 � $TIT1d ��� 7Td�7T� 7TP7T55V6�5V75V85V95W0 5W>W�A7URWQ7UfWU1pW1zW1�W1�W� 6P!SBN_CmF�!�0$!�J� ; 
2�1_CM�NT�$FLAsGS]�CHE"{$Nb_OPT�2�p�(CELLS�ETUP  �`�0HO�0 PR�Z1%{cMACRO��bREPR�hD0D�+t@��b{�eHM� MN�B
1�U�TOB U��0 9DEV�IC4STI�0� � P@13��`BQdf"�VAL�#ISP_�UNI�#p_DOxv7IyFR_F�@�K%D13�;A�c�C�_WA?t�a�zOF�F_@N�DEL��xLF0q�A�qrc?q�p�C?�`ıA�E�C#�s�ATB<�t�d�MO� �sOE � [M�s���2�REV�B3ILF��1XI� %��R  � O�D}`j�$NO`M�+��b�x�/�"u�� �����!X�@Dd p{ E RD_Eb�~�$FSSB�&~W`KBD_SE2u�AG� G�2 "_��B�� V�t:5`�ׁQC ��a_E�Du � � �C2��`S�p�4%y$l �t$OP�@rQB�qy�_OK���0, P_C� y��dxh�U �`LACI�!��a���� FqCOsMM� �0$D���ϑ�@�pX��OR BIGALLOW�G (KD2�2�@VAR5�d!�AB e`�BL[@S � ,�KJqM�H`S�pZ@M�_O]z���C�Fd X�0GR�@��M�NFL�I���;@UIRE�84�"� SWIT�=$/0_No`S�"C�Fd0M� �#PEED��!�P%`���p3`J3tV�&$E�..p`L��ELBOF� �m�@�m�p/0��CP�� F�B����1��r�@1J1E_y_T>!Բ�`��g����G� �0WARNMxp�d�%`��V`NST� CORz-rFLTR�/TRAT T�`� $ACCqM�� |R�r$ORI�l.&ӧRT�SFg���CHGV0I��p�T��PA�I�{�T�!��� � �#@a����HDR�B��2�BJP; �C��3�4�U5�6�7�8��9>���x@�2 ]@� TRQ��$%fh��ր����_U�������Oc <�� ����Ȩ3�2��L�LECM�-�MULTIV4�"$��A
2>q�CHILD>�
1���z@T_1b ; 4� STY2�b4�=@�)24����@�� |9$��T�A�I`�E��eT�O���E��EXT����ᗑ�B��22Q�0>��@��01b.'��B ��A�K�  �"K�/%�a��@R���?s!>�O�!M���;A�֗�M�� 	��  =�I�" �L�0[�� R�pA��$JOBB������`���IGI�# d Ӏ����R�-'r��A�ҧ��_M��b$� tӀFL6�BN9G�A��TBA� ϑ �!��
/1�À�0���R0�P/p ����%�|��Bq@4W�
2JW�_RH�ECZJZ�_zJ?�D/5C�	�ӧ��@�����Rd&� !����ǯ�rGӨg@�NHANC��$LG/��a2qӐ� ـ@�B�A�p� ���aR�`�>$x��?#DB�f?#RA�c?#AZt@��(.�����`FCT�����_F࠳`�S	M��!I�+lA�%`  �` ���$/�/�� ��[�a��M�0\�ؿ`��أHK��AEPs@͐�!�"W��N� �S'�I��' � . II��2�(>p�STD_C�t�1\Q��USTڒU�)#�0U[�%?I-O1��� _Up�q��* \��=�AO�RzsBp;�]��`O,6  RSY�G�0�q >EUp��H`G�� {@]��DBPXWORK��+��$SKP�_�p��DB�TR>�p , �=�` ����Z m�OD3��a _C"�;b�C� �G�PL:c�a�tőS�D��G�Bb���؎P�.� )DBd�!�-|B APR���
�@Ja3��. p/�u����� �LUY!/b_tS��0�_��/�PC�1�_�T�ENEG�]� 2��_�S6PRE.��R3�H $C��7.$Lc/$USނ�z )kINE�7A_D1%�ROyp��ŀ����qbc7 T@zfP�A���RETUR�Nxb�MMR"U���I�CRG`EWM��0�SIGNZ�A� ���e� 0{$P'�1$P� &m�2�`��`tm�pDIp �'�Bd.a|	r�GO_AW ����0ؑB1m@CYSd�(�CYI�4��B�`1wsqu�|t2vz2�vN�}��E]s�DEVIS` 5� P $��RB���I�wPk��vIG_BY���p�TQ޻tHNDG�Q6� H4��1�w��$DSBLC��O��v�G@�Ǝ@_qL��70/�F@]�d�FB���FERa8����t]s��
�8> i�T1?���MCS솀�FD ���
[2H� W��EE���p%F��ŻtSLAd��09  ��INP�^��]�`�]q��:P +8�S��0x�`^���^���FI�2�������A	A9Wl���NTV�㜒�V~���SKI�#T�E����a���T1J�_�#;2_�PD�SA�F�T�_SV�EOXCLU�῰�%D6@Ll �Yք��3�HI_V
0\2PPLY�@0«�G������_ML%��pVORFY_�C��M��gIOC�UC_� ����O�p��LS(�`V�&T4�A1��s	���@PdE&�gp�AU��NFT�u��upZ��pm�ACHD��O���^���AFC C	Pl��TD�4P~�� N�� ;�P@T��|�0,@ ��I�r��N��=� <Y���T��?� ���{��SGN��=;
$ �`�a>aR0I�3�g@� _BM�_B]�ANNUN�P~��ÅuC.@�`/�ɢ�� �ʬ���2EFC@I�R>�p�$F���4OT�`{�&TD�(RQ<�j#QmJ�Mb�NI�R!?��4һ6�A��R��DAYCLOAD��tT-�'S5#Q�EFF_AXI��%@�PQO3O�йS��@_RTRQ��A� D1�	`��Q,@ ��EVp�Ӓ����@�0}�0��{��MuP�E{� BV������$s��DUt�`����BCAB��C���PNS"�+0ID�WR���V!� �V�wV_���V ��DI� �4D� �1$V�`SEm�T Qj}�'���D�f^E_n�$�VE� � SW���[�a�����A��O�H��)�PP��%�I	R�1Bu@p�&�� �b����]�w3W�O � W��vM���C�0��cp���RQDWF�MS�w0��AX,���$�LIFE�@����-Q��N������C�o���CB0LqN0]a���OV0sHEQ�SUP�T����@_oS�1�_��Gq�Z�
W��
B1��#��@�k2X�Z_ LQY2�C"9`T_@``��N����*��J�! >�_� ��xF� �4E `�p�CACH,�\�]SCIZ(T ���bN�oUFFI� �� �@(T��'S6#Q�B�Mp0�F 8��K�EYIMAG�cTM,aV#��a�^�hB>1�OCVIE�a�G�2� L��H���?�� 	��D� PH����ST'�! C"D�K$PK$-�K$��>K EMAILK�u`x[��0��FAUL�R�I�2sc�C� COUȳ0iA�0T`�1JO< $�#�S�vm�ITW�BUFp���p�t�0�0n B�$�tC�����"�3� SAV-5�"����H7@@��P44�
`��N�_� 5LЉ9OTgb+���P�P�:����7AXC����XX� T�a3_G��
m@�YN_N� K <�\�D�uPb�M�M�8�H TL�F~`Y$�`��DIزE�@H`�aLY���G1��&G�Da:AF����baM�`A�#�3C_^`�`Knd�@^�DQ�R��E�(AD�SP�BPC�KI�M:3�C�A��A��U`�Gd meڠ� IP��0C7�3�DTH��d�B��Taa�CHSEC��CBSC	�"�PV����Z�P�3�Tp��NVk�G�S�T�F� 	F���0d�C5@�1a�SC���u�CMER|��QFBCMP��v~@ET;� N�FU� DU� ́�`���CD�IYP�0�#�m��`NOu�=�O����pzbL�xds�P�zbC"��e
��2��!uc�0� PH *�aL��_c�q�1 f��,�'��dD��f"р�f-��f���f��f7
�i8�i9�j���hzU1z1z1(z15zU1Bz1Oz1\z1iz�2wz2{z2z2�(z25z2Bz2Oz2�\z2iz3wz3z3T{z3(z35z3BzU3Oz3\z3iz4wrN�EXT��=�QB \h@%@�e@C��e��0FDR��RT� VW��2��\�R��REM��FqN��OVM�C��A��oTROV��DT806КMXߜIN��: �Ϛ��IND���
�F@�0@G�1d�ِ�9 ��D��ِRI�V԰&��GEAR��AIO��K��$�N 5@��������� %�Z_MCM� ����Fe UR3bS y,�a1? 9 �P?���?�E,����1`v��T���P�1��R�I^e���#ETUP?2_ U -��##TDGP0��$Ti��pZ�T�qa�"BACBGV TD��"eD)_J�%�ýc0@ѰIFI�:�0@`�`�Ь�PT���LUI6$Wc �� (� URt� 1@�2MA�P� �����I��$(�Sܰ?5x4�Jb@CO|0�3�VRT$���x$S�HO�ѱ��#ASS�jP�1(IPQ�BG_ ����s��s��(s��5sFORC�"7�籯DATA��X�"F�Uס1:B��2:AL�OG���Y |�*�NAV�0��(�X����S�"&�$VISI[�.BS�C�4SE�t�7�V*B�Or���Bò��A�Z�$PO,�I�E��FMR2>s�Z ��i` f⁑s@�օ�������Pǖ� �堒_wqX����IT_ֱSd��M�E�j�|�DGCLF�;�DGDYd�LD��H�5
?�ѡM�cp8#[��� �T�FS�07$\ �P2���sC�0$E#X_������1�0�P�E��3�5��G��Q��] ��0bS�W5O��DEBU1G��]�GRc���U�SBKU`O1n�p  PO�Р��t�"`G�t�Ms�L�OO�3��SM�E�<2|��& _E �^ ��TER�M��_��� ORI�SA��`��cp�SM_`@]���a������� b��~�UP"c�� -�D�^((���f _>�Gk
}�/ELTO�!>B�PFIGf?AנS�`|b`$UFRfB${`�� Ne�3OT��PTAiP����NSTT@PATx^Qi�PTHJ&a�L`E9 d2U`�AR�TU0�� U1�">AR�ELAc1SHFTPPR?A3__�R/`�Ic ) $8�b�.႐S�S�2SHI�d+�U�b O1AYLO.P�1 A��j�p���e[PERV p �$��T@A��0Ȱ+%��ȰRC��e�ASYM3A�e?AWJ�$� �E$�/[)�OaU$T@ A3���&IPS��Q�O5RT@M��/�����d��t��� �1�6�HOs���e �˶s�i`OC�|��$OP^��A�cv���a�i@���R0R�S"OU,�Se�R�5�m8K��e$PWRf]�IM�5"R_H3`(*� ?AUD$�FkSVoc1SDfH��$HdE!@AD+DRC�H��G7A�,A%A"�p@F��ag H2�S�PFѝ�dE��0dEsdE(sSE��HӶ�`HSY`MN�hW�@0��"QebaOL/SW�{0R�\f���ACRO����ND_C/Szb��4�QOROUP�S2_��
Ғ�11�q��:S� DY3 DY��EXpDY(p�DY����AC���SAGVED?W�SOUG�C���i $��@0_�D)���j«BPRM�_
�~�HTTPu_z`H�aj (;`�OBJB�%B��$�C�LE�0a�`k� � 4��6�_�T��XbS0�3���KRL�9HITC#OU����G�LS�j0�Xbb�$�f�j0ʷk0S�S���dJQUER�Y_FLA�C_ _�WEBSOCI���HWcq�+�l_@>� INCPU�R*�Ovma��K�0pzD/q��D/qǂ�IOL]N��m 82�R���i�$SL��$�INPUT_���$�0~xPy� m�ZpSL�P+�nep�{�u�tB#�uB"NAI�O�PF_AS��oF��$��B��qN�Y��2��ksM�ts�HYB�5���A�pwUOP��p `�p S�C���%���,�}��0P�3�0s���,�����>�IP_ME\��7q X�pIP,@�R�ւ_NP��`*�`G2B��O��BSP���P���BG�Q�-�9M<!�r l ��TA�3`As�TI����%� ��_�OPS6^�BU��ID�Ўb s���x0��;a-���� s�r?�r�S��p�NҘ��ӕ�IRC�A_CN� tk �Ji�pCY�@EA��C��q��3�1�#��@z"���!DA�Y_����NTVA�����u��r#��u�S3CA�u�CLO᎑"j����@��u��ڔX$��N_R0Cβ򐎒c�6�v�r��^3 %���'b�����Pi���? 2u �p.�����w��\�'b\�L�AB�z��Ѐ�UN�Iбn�	 ITYl�.�0EL�R; G����x�r�R_URLnЀ$A�AEN|��k�*��0�CT�AT_�U#� �Jp��y�р$�_%E�pR�k�.��AS��q8�J��aC�FL��K��P
|W�r�
�UJR�%z �J`F��(�����D£$J7,S%�J8��7&�h�$����7���8�ɭ�oAPHI�Q��z��D��J7J8"��L_KE�� o �KQpLMܑ� { <٠XR��p$p�WATCH�_VA�A�ű#fF'IEL�"Cy�2�&��| 
��V�G-1���CTܰ�������LGɳ}� �!�LG_SIZ�Rdv��հ����p��FD��I���ة����� ������d3��V��V� �pV��V���V�K!G�:� _� _CM�������F�!������r�4(�Ѡ�р�������p��� �I���
�����������RySU�  (��SLN���"~_��`DE��E�r!�s����S��0L���DAU��EA�PQp44��Ʋ�GH52X��pBO�OYA� C�ʀIT�c��� �sRE4�SCR���|c�D�PKr,QMARGI�q�;�v��S4e�d�qS8c�rWpC�q���JGM��MNCH���qFN�(ҞK����	UF����FWD�H]LSTP�
V��������RS?H� ��C�~"�� w�U�Q�v�����G�	PPO�"2�� �v�	EX�TUI�I;���;�8bZ#�Z#� ���R��P#� #N�A�3ANA�rA1��AI���D�� �DCSf�lC�#zC*�"O�(O�'SK�2r�(S�(ZIGN���������4��$DEA|LL"�Xp�q����Ѐ�м�T��$@�׳�r
���AA���۠lp*s�A���S1�52�53��1.�"� �Ђ �Jk�0�$�u�t����Q�e���:FST�e�R��Y�B\A /�$EkFCkK����PzF�F{�$�у Lp#�n�8����Co`���d�P�D�5#_ �X�Np�Q��$ �Sp�MCt��{ �J`CLDPe�> �TRQLI��"�PY>TFL%�iR�QrSb��D��rWpLDrU\TrUORG(�v�R~��RESERV2t��T>s�TIr /Sv�� � 	[UvMTFrUSVd�PP^�	�Q�+d3fRCLMC�Ad�_�_SiTp3al0M�DBG�qͰ�?��$DEBUGMA�S&�_�P���UuT�� |�E����PF�RQV�� � ���HRS_RU��q�A'�A5��FgREQ����$� ��OVERt���tF��P�EFI��C%�A(��a���c��T� \�q��s$U@%�?`���PS�0C�	sC ��BcN��sScUݐ�a�?( 	{�MI;SCuŊ d}�AkRQA�	�TBN ƕ� �m!�AX� �-��.�EXCE�S벿��rM��̱�½��r �Q�rSC>@ � H"�	�_S��8���,�>��P�Kɴ��r��N �eB�_��FLIC�DB� QUIRE�MEO��O�pv�aL�@Mȵ� P��E�h���AbZ�ND��q�ހ�{�r��؄�D|���INAUT4���RSM����+0N�$bn�j�PSTL�̱� 4٠LOCfFRI��EEX��ANG�"�q�aOD-A�e��p|����MF���Cv7I�B�A �Eq�o�fSUP��FxpFX;�IGG> � �`�C n�(�C��Da�br\B ��^@ɨ^@ئ���P��7�qTIvл�'��0�IN�b� t9�M	D6���)D�� O�Xa�L�H���O�DIA��P�>�WiO��1�
O�D��)/�t�)`ހ�� m�CU��V ��#`�q/�\_�`y�� ���CC��`rr�� �P �J���P��KE�^����-$B+p��@ND�2ZbZ�P�2_TX�DXTRA�#|�lbM�E�LO��ހ�k�L��� ��u�ǲ��ƪ�m�RR2�u�O� .����A0a� d$CALI��o�G�!��2�0RsIN����<$R���SW0_d,�lcABCJ�D_Jb����p�C�_J3W�
Q�1#SP�Т��pPQ�xݡ3w�̱�@�p��J�lc���R(aOu1IM<l`�rCSKP_Z��H���#��J���rQ���������_AZ/b��I�ELZ1��ZaOCMP��q�q��cRT�at��1��Ќ���1���{ ��Z���SMGY'�zdJ�GPSCLN�
�SPH_0�p7��㓰z�p��RTER+В��� ��_� )Q�6@A\ SC�r'�DI�_���23U��DFڬ0H�LWN�VE�LPQIN�Bf q�_�BL� �ry��ѳqJ�i�~�����MECH�2lb%�IN
�q��!�ǲ��]�q���@_�p �����/���0�􆂛��?��0D�HN�~�����0$aV������{!$��X'qrA�$O1����u�H �$B�ELZ��g�_ACCE� �la� OIRC_(��a�P�NT�q;C$PSN�CRL�0��XS ���?�� �G��	D�3�ؠQ�_�1�lIO"u�p�_M�GsDDl(�rFW3P(�����}�DE�PPABN6�RO��EE_�1 �PP��1�a����0?$USE_���#]P+pCTR�$Y��~ .a �AYN�pA m 6&��f�6!M�aұ��"fOk�
c$INC�������'��.�ENC�L��r����� INCBI0��%)���NTi��NT23_L�r�#CLO]�r09pI\� �6R���p���0���C���&MOSI�q��߰O!s�rPERCH  ��7q� y7��3�2zd�@o�g� %&N��AC�5L$�ӻ����%��8:F36TRK��AAY���3��HACWE�LC�z暁�"�`MOM}"����P̰�����cC���DU���DS_BCKLSH_CC�E�`X6 8p>#�s�C�"ZM!�CLALM�$�a�@ 5UCHK���Z�GLRTY��A��$���Q'�_f�M4_U	M�c�VC�cz��SnpLMTt�_Lj b�Tv��WE�]�P�[ �P��U��нc�2 d&�8PC�1�8H��&�p�UCMC��z~CN_	�N��f��SF��9V "��'��TaC�eXhCAT�^SHf�	�~�&yQ��A�&����ɗ�mP�A�T�"_P�UrC_ ����OFm0��_CqtbU�JGJ�d�esW�OG|rg�TORQU  ��K3hI��c2��r_W�EHD��m�tP^�ud�uI�{I
�IdF0��q��I���vVC� 0����j��1p�n��0�v�JRaKp�������DB���M����M��_DL^�2GRV�t�^�dՁH_��Ӄ�"�COS/�|�/�LN��R�s�Y�^ T���@T�&���~�D�ЅZM�c6ՁMY[�Θ;�I�|C��THET0#5NK23d�X\�[CB�CBXC��AS�C�&�Q�^Q���SB^o�)�GT	S���C{�Kq��:sx�祪��$DU_P@�7ʢ��٧��Q�1Y_4cqNE��AKoT��-�< �A��:�C�!�,�,�LPH/���%�Ss���~� �������������:�EV\�VQ�N t�V��UV��V��V��V��VȻVֹH\�u�{�Ps��a�Ȑ�H��H��UH��HȻHֹOM��O\�O�r�O��O���O��O��O��O
ȻO��F�>���~����O�SPBALA�NCE_ޑ��LE6��H_�SP��o����~��ҍ�PFUL�C����⍕��1=���UTO_ZPbU�T1T2^�2N AQ�� ~���A���(���AT	@OA�>�pINSEG�<1�REV��<0�!DI�F2E	1���?�1�%@OB��%Q���G�2�p� LQ݄LCHgWAR�%"ABAq�E��<0ސU!���SXUAPdt�3�?S��� 
u��q��%ROBm0CRC��ib���C�_]rT �� x $W�EIGHR p$�M���tpIR!0IF�
!�LAGC""bS�C"��C"BIL)O1D�@?0ST� P��%P p| �`��
����
� �D!]q�  2�J4DEKBULXɠOMMY9���N+s��p$D�1�$� op � _ �DO_� A��� <��rh��D!�0�BB: N�#_�!0D  _O2P _�� %�PT� ��!�QT��� TI�CK-�T1� %j�@sNm0M�	m0R�@D!=�=�� _PROMPR#E/�? $IR�pB!phP��0"MAIڀh}!T"�_# ����^AV R�COD�wFUJ ID_��0'%�����G_SwUFF&� 49!��DO����< �GR#=�e$ �q$=�|%=�%�qe$��� ���H�_F�Iv9�#ORDfB ��36b��"B!� $ZDT�.%"@_��4 =*��L_NAs|52�DEF_IE8 52�Q4�I�S�0}3��5�IS��` ���3�O4�a"�4�abSDQ��B��4wD�pO�� LOCKE+q_#��0��1e"_ UMd%52 e$}3e$�5e$�2q"gC p%`3q$�4q"Q�F�1 |#H�^q|%52|%}3|#�GUa(8P�4H��1�� WFHEU<C?���TE0Q�ߣ LO�MB__RzW0V�IS=�ITYA�oqOCA_FRIN�S�SI�1�Q�!Rp�W{�W3��W�XW�[倩V��_i�!EAS�"�q��Tp@��V4�Y5��Y6ORMULwA_I+q�G%7_� h �7�COEFF_OW���dW��GqS �CA���_�GR� � �G $<@��
XGTM/G't<E]DCA|ER��T%D$4� 7�  G�LL�$@�S/�_SV�4�x�$hV� ����d� �{ rSETU�3MEA�D b� _|�"�� � �p�� � �` �� ��A�:2sA0AD�b�Q�";��@A�1@G�����REC�!�� M�SK_��s� �P��1_USER�z�j���,𾔙�z�VEL>���,�����=�I0���MT8C�FG���  �u��Oc�NORE��� ��-��� 4 �s^�d�XYZ�#����d���_ERR��! ��ep6 �c\��}��Ҁ� BUFoINDX1�  W�wMORt� H��CU\�d��1xӃ���!$������10��a���G�r� � $S�I�`�P �ᝀVOx
����OBJE��ADJU����AY9p���DJ�O�U� 5���C!�"=��T��y���x��DIR}��������⎴�DYNb�b��T�R�5�R�QHB 4���OPWOR� ��,� SYSB9U*�2�SOP��$�q�U���P<@߂4�PA���6�_�2�+OPz U4�(��xt�e�IMAGo�1��q�SIM���IN`\���RGO�VRD��%���g�P i��������@ C׵d��L:@BY��� �PMGC_E0��N*�M±�1��p��sSL���� ���OVSL��S:RD#EX�1�0K�2c���a_��cǬ ��cì  mÂ�}Ȫ��C��70����Ƿ�_ZER� �*��s��� @h"���~�O/ RI���
��������T��'�L�����T`�W ATUS�p�C#_T����O�B+pYրB���3�.�0��� D�e�N�LҾ��`M��!��o��XES� ��һ҆��ò�����R�UP:��0�1PX��y�b��3ǂ� ��PG텳��$SUBA�~��AA��JMPWAIT��r�Y�LOW/�^�' CVF�vc�\�R���q�CC��R���i��IGNR_{PL�DBTBW P�1d�BW ����U*��IGL��I�c�TNLN����R�֡5B�PN�E�PE�ED��T�HADO!WW b���ES�M��b�+�P0SPD��� L��Ar�Q0m�/��{�UN �y���R�м�LY0��Kѓ�^*�H_PK����?RETRIE��bi�'����FI�Ƕ �:����� �2���DBGLV~��LOGSIZ���1KTy�U�s2D�8� �_TX�EMB�`Cn���X ARR|.R+�CHECK��N1��P��p�c������LE�4pP�A#@T��C�O��P4��p�bAR%"���#�1'�O� 0��`ATT���x�%X 0��1��UX�����PL,  $���/QSWITCH�T��aW�AS����SLLBp��� $BAv�D
C2�BAM�������J5L����6�|_KNOWh����U=�AD���`x�D��)PAYGLOA��@%#_���.'�.'Z+#L�AA��q�0LCL_ʐ !�pg"�Ӂt$*˲�&F�)Cgpb*(�e$�`Ib(Ripb'${�~$B7`ʑJ���!�_Jl!��֑ANDz�U�
4l"�!(�"a�PL�AL_ ��`x�ѐ����PC�>�D*#E=��J3�036� T�`PDcCK�22�CO�p�_ALPHC3�3BaEБsaC?U< ��b|��� � �.�$/D_1+*2U$D�pAR��H�5FC^�TIA41I51I6>�MOM��=C]C�JC]CWC�Bp�AD�=C�FJC�FWCPUB�RbD�EJC�EWB'��@30ʑq�  �� MO"L� ��T���� e$PI����3��0'P&Y��J)&YI2[I@[INS�DS�V�V�ޠ2������1�HIGo1�q�j��Vj� q�����V�S�X���Y<��q�SAMP�Я��:d�W;cq�3 �piaʐS�Œxd� �fj��0�i@Œߠ䢐:@�e/0��H��cIN�l/0c�h�k�dq���jx�d{2{GAM�M�eSU�A�$G#ET�R��3�D�4҂;
$60IBR���]IL�$HI:�_��H��Œ�vEѐ�xA�~�p�vLW�}�v�|�y@��v�2�V�51C��GCHKİ��q�x>I_`�ޔ.2�8.1��e|�uCޔ�F{�33 ��$e8 1���I�RCH_5D����RNs�8���LE���R����8�Ѐ��MSWFLܡ��ASCR�100{�. xd39]��g�ʐ=@�iq�j���PI�3AVMETHO��æ��妒AX$���X4�p�ERI���:d3fsR�� 5	D�Q�0FWt;ac��c�(�L�;a=�OOPa֑S��a֑'APP��F� 0W�x�c��cRT��2�O0j�0�������DR 1�%��D��ѪNP�ѢRA� MG�vOSV	Q�P; �CURC��GRO<7���S_SA�ܴ,5���NO�0C���� �45��t�?6/H/TX�����zP��UϸCDOi�A�rdyes��e�X ��W��X3�/��k#����D�T� � ���YL$S�!�g���S�"6A9��K����!�����!_�C����M_Wd���C�����?�M���ˇ ��21~�L�T�K��r PM&�R� ��}�R��WE�S$��L3X!EШ4Cү4@CҶ4C�W4���pN�P�sf��/0X��O�3�.1Z�� P{�T� ���M��z�w����������4@����� ��� P�1_Z� |v1��5�]I��JC�� WC5�6J���PJuu(Ms��ſ�Y s��P��PMON_�QU?` � 8�� QCOU��Q�TH_�HO~�:�H�YSES�:�U�E%�+�� OX� � ��P#ПuV�RU�N_TO��o�O��R
P� P! ��Cx����INDE�ROGRA��J��}2C�NE_NO��ƃ�IT�A��g�IN;FO��� b�������  �����{ (SLEQ�V`"�U" ��A�OSU���� 4� EN�ABqҁ�PTIOyN
�ERVE�Rp~�Q�VGCF_� @.�J �.1��+��pR��|=�T_EDIT��'� �R���K�A�S5�qE�pNU�AUTQ�	COPAY�A�P*�Q]�M�q�N48M�PRUT�R ;N� OUC��Q$G��?�R�GADJ��� hv0X_��I���п�пW�P�����S��rN0_CY�Cq��RGNSr[�s�=�LGOZ���PNYQ_FRE�Q�BW�`�VP!SIZn[�LAœG!�8XC�`�UCRE�p��f[�IF@Q��NACa�%�$_GœST�ATUv�œy�MA�ILAb�1�!
�5�L�AST�!�1"$EL;EM_� �\�iFEASIl3�nb g�Z�2��>�96���`�pI����G"�Q=� �L�n2ABU�0E��r�PV�!�6BAS�2��5�r�AU�P�PJ��$�1�7RM�@R h3Ł���3���P�r�!ƺ4 ��$"S��~�	E2 2� �c���d+F�2*G�2�"Э`���2VGW�DCOU����r�"$P �z@�)GRID���U�BARS�WTY�m "OTO�����+ t�_�$!��B�DO��\� � 9����POR���C\���CSRV� )T6VDIS�T_�P4P�FT�PPW�PPW4NY5*NY6NY7NY82Q�Fbr_�r�$VALU�3(�+4)0��}F[�� !h�^����C�!%���A�N'��R�!��T")1TOTAL_�$l06b�PW=#I�AKdREGGENIj^b��X�8`��=�� f �TR�3�"Ia_S+��g^`��AV���b��2E�#� �?�(2�� cV_�H�@DA ��`pS�_YY���a&S8�A�R �2� �IG_SE6�`R�%�_���dC_�F$C�Mm�f�wrDEh�?p�rI]�ZvsPsq!z�F��HANC&�O� pAj�"d#qINT1P��yF}���MASK��0OVR��� �<�0�!Ł�Gy�,�Q�E��d�OJ6�k�F�P�SLGHp�Q� \ 1�b%Z�$�3`� qS���$�qUY�`y����c��ZQU d��w�TE��@� (�aJV�Q�q#OIL_Mp$�Vt2����TQ ����0�C���VB�CP�P�_�J�Z�Mq�V1Vp�V1~�2��2~�U3��3~�4��4~��� ��<�����IN�VIB0�J�7�T�>�2:�2F�3:�3F�4:�4F���Y� r�U��gP
�tP���'��PL� TOR$��IN��u�5�����T $MgC_FC�X���LC�B��u)`M��I�s*�rC ��)�r���KEEP_HNADD#�!e��0o�	C�ѳ����A$�����O�d�>"��`��\�w��REM������!�Bµٱ޸U�$e���HPWD  �e�SBM�q�@COLLAB"��P��4'a�" IT' ���INO)�FCAL�h�
���� ,��F�Lnб1$SYNT���M��Ccr��`�UP_DLY���r�DELA���!�"�Y �AD �.�Q�SKIPG�� Ą
P��O��˂K���P_����Ƕ���� �#ٖ#�gP"�tP"� �P"ڎP"ڛP"ڨP"�=9��J2R ���dX�0TJ#���� )1�Ѭa�����a� �RDCaw�� �� R��R�!�=��-DRGE� W3�{BFLG�0��S9W{	-DSPC��!�UM_����2TH�2NuA��� ?1� ����A>[ � D���x<]�02_PC����S���1Q L10_�Co"�ѩ��q ���JPٰ7��6K�@+��� �.�NE����N���b\r�3�k����p����DE�SIG��JEVL1b��1��k��10ٰ�_DS�K���ڧ�FC11��� �lV�������iI�AT����AS'J N�$	C�
���HGOME4����2������� 2D +,��3���gy@���� ��4�����,> )����5���as�����V6�����//&/8/P7���[/m//�/�/�/S x��8����/`�/�/? ?2? ���S)����  @�1��s`Y�V۰E�D� T���4,f�3�IO��
II�0XrOe�_OPE.C&b�3��POWE��# �0������&d� �}�eB$DSB��GNAr�%c���C��t��S232N�5� ��Z5���׀ICEUS/cS�PE���QPARI9Tq$aOPBQ��RoFLOWApTR�041b�UJsCU�@6���QUXT�q�Q�pEORFAC�DʰU `�VSCH�Q� tV��_�@kpc�3$�`�`OM*p���A>�#�p%�UPD�<����aPT�0|uE�XЙX|S!%�FA�?��rj�r�a � ���`;b K�AEL$� ��U��]B��a  2� ��S���0�	� ��${�����GRO��`*dT�(p6fD;SPBfJOG�`�C����AZ�N�������"VK�P_MIR�^a~d�MT3��cA�P%����`}t��S�p�`R��
��eBR�KHUQ�V��AXI�1  �bc�r-b��q9�7e�`BSOC�6f۰N2uDUMM�Y16O�$SV&��DE3A�CF�wK�e0�D�pcOR{ws0N�p|vFp�w[`�OV^eSF�zRU�N�s�rF�vQ�cU�FRA�zTOTLcCH�����OVlt[�[`WP�7�[c���r�?p��_�p� @>h�TINVEG@n1�OFS\�C�P�WD�q��q>qf2�eXp�TRr��1a�E_�FD�aMB_CW���B��B�*��ałˁ?�epV9Q��P�&��írGƇ�hAM��c��VP�F�!�_M`݀R_�CS�T$�����Q�3T$HBKX�Q�fm�IO�5|�&A��PPAp�����ଔ��,�&BS�DVC_DBъ0ސ�Q�B ސ7�Q������F���3��L�E���+P�`lqqU�3P`FCAB�Ѐ�2~㷀8û` ���O��UX�fSUBCP�[�-��/���P/Ѯ�ރ�bB��$HW_C��	P/ш���?�q0#��P��$UP�t	��A�TTRIh��h`C3YC��g�CAB��c�FLTR_2_FAI�3�IH��F��Ptk�CHK�_SCT6�cF_�F_�����FS�A��CH�A�}�ֱ�RղRSD���Aq�S�A&@�_T�}�.���PE)M�0��MsTò/���Pò��K�DIA�G�URAILAC4듑�M`LO"p��<Hv_�$PSNb�2� ��L��PRߐS�}�I���Cёf�	�E�FUN��*QRIN1�}�|0^���Q&�S_;`��X�����0f���P�f�CBL���.�A'�#�*�#؃DAp��h�.�'�L�DyP`p����Ca�����TI�°���P�$CE_RIA�a�BAF��P�AX��~���T2}�C�S��؁OI����DF�_L�0�r�Q�PLM��F^�HRDYO,�af�RG��H���a�|0p�/�MULSE������Qp�$J�xzJ�r�w�{FAN�_ALMp���WR=N��HARD�0�VZ0P]R�2���A���e_��fAU�R�ȴRTO_SBR &E�O`#��ӓ��;�_MPINFQ���N��Y�REG�6NQV�Pf3�fDA@N��sFL��R�$M�� ��`S����P�����CMѐNF-��1�����h��A��0$Δ1$Y oQ�b�Q�0�� ���cEGI@+c`p+A1R=`CHu25Rr:�T��eAXEEgRO�BBjREDBfWRd,� q_�$sSY�`�ep�S�WRI,�>�STr@CcP�p�pE��0G6�Rr��;`B� R��7\��2�OTOi��0��ARYBc4~�2�̳2t`FI�`�c$�LINK�GTH�S�PT_�R�rF8Rr|XYZ�R:�9�OFFZ�S){o8B@`����/��@�P�FI@1�����CXt��Zd_J�A�R�r`����30Rr�@�*!dm�b"CFA�eDUn�rHu3����TUR��!X�ӛ%BI�X� `�J'FL|�a�8 � ԝ�	3ʡg� +1��0Kg`M�d�&�Qs�����°�pSOR�Q&�Oa�P(���`O � �1ɐj4��Ma��~4'OVE�1MIPk1 ��5�5�6_Q�70c��7��4ANڡV �1���1�`�0�k1 �5�1�7(E(E�3OaSERla�	��E,�H�P��fDAA�P����!�@o�l�o�AX /��Ro�2��U�EQ� �I{��I���JN �J��J$�J��J��J1 [ �F/��I/��I/��I /��I/�Y/�Y/�(Y�/�8Y/�HYeQYYDEBUڣ$����U�	ao�wABo�m��qr3Vb�٢ 
$b �LeʡXgQqXg�� XgNXgXg$Xg��Xg���g ��U�L�AB�J5֠�G�RO[�J"��K�B_/�MF��s� �v�5qK51u�=vAND 0��[DL��^A�zw K���� �x1ѝxN��NT��#��pVEL5��4�qm��x9���NA��m��$���ASS  �����* *  ��_�SI@���#��)�I�Y�n��(�AAVM���K 2 T�� 0 � �5�����\���� ��	݀΍�* U��ߏ��!�͌@�L�܁R��������e�BS�1  �16�� <u����
��.� @�R�d�v��������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ� �߲��������߱��p�MAX/� ����ʓ  d�IN��*��PRE_EXE;�g�J�!43���T�e�IOCNV,�"<� �&�P��a �;�Ɨ��IO_�� �1r�P $b��`���V���U�?��� ��$�6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�o(:L^ p�������  ��$�6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z��������ԟ����LA�RMRECOV �~�!�J���LM_DG ����� �LM_IF ��+��ߥ���ɯۯ�骓���0�B�S�, 
 S�|���@�����ƿؿ�$�� ���1��U�g�yϋ�����NGTOL � ~� 	 A�   �����PPINFO Z� Y��*�<�N�!�  f�P�~�?�m� �ߑ��ߵ������%��5�[����χ�� �����������)��;�M�_�m�PPLI�CATION ?}���g��Handl�ingTool ��� 
V9.1�0P/30��j�?
88340�����F0����1028��������7DF�1��j���None�j�FRAj� �6w�_ACoTIVE�  �����  �UTOMOD� ^��Ê�CHGAPONL�� �OUPL�ED 1��� �
 2�CU�REQ 1	�� � T<<<	�����@��<�����Hk�HTTHKY�A�o�� �////�/S/e/w/ �/�/�/�/�/�/�/? ?+?�?O?a?s?�?�? �?�?�?�?�?OO'O �OKO]OoO�O�O�O�O �O�O�O�O_#_}_G_ Y_k_�_�_�_�_�_�_ �_�_ooyoCoUogo �o�o�o�o�o�o�o�o 	u?Qc�� �������� q�;�M�_�}������� ��ˏݏ���m�7� I�[�y��������ǟ ٟ����i�3�E�W� u�{�������ïկ� ���e�/�A�S�q�w���NTO����DO_CLEAN�|��NM  �� <_�qσϕ����BDSPDRY�RϊHI� ;�@ L��%�7�I�[�m�߀�ߣߵ������߇MAX~�������	��X���PL�UGG� ���P�RC��B9�=�����c�Oh�����SEGF� K������ 9�K��%�7�I�[�����LAP������ ��������	-?�Qcu��TOT�AL+�T��USE+NU��� ޸���NRGDISPWMMC��0�C��&�@@���O�������_STRI�NG 1
�
��M� S�
�
^_ITEM1h  n���� ����//&/8/ J/\/n/�/�/�/�/�/��/I/O S�IGNALb�Tryout M�odeiInp�0Simulat{edmOut,<OVERR��� = 100lIn cycl 5�mProg A�bor63m4S�tatusk	H�eartbeat�gMH Fauyl�7�3Aler�9 �/�?�?�?O#O5OGO8YOkO}O ��d ��v�O�O�O�O__ (_:_L_^_p_�_�_�_��_�_�_�_ oo�OWOR��dJa�O$oro �o�o�o�o�o�o�o &8J\n��8���~POb�1 �pbk��#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g��rDEV�~������ ˟ݟ���%�7�I� [�m��������ǯٯ�����PALT �M6�bo�^�p����� ����ʿܿ� ��$� 6�H�Z�l�~ϐϢ�$�GRI�d��N��� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F���� R�M~� ��X��������� � �$�6�H�Z�l�~��������������l�PREG:�# ����J\ n������� �"4FXj|���-�$ARG_�J`D ?	������ � 	$�&	+[�]���')��SBN_CONGFIG� �$1#2�=!!CII_S?AVE  �$F!�9#�TCELLSETUP ��%  OME_I�O�-�,%MOV�_H� �/�/REP����/�UTOBA�CKv!�@"�FRA:\ ��/F '`�0�C8� T;? � 23/0�7/18 17:_50:04(��?�?�?�?4<�� O6OHOZOlO~O�O�$O�O�O�O�O__ �O<_N_`_r_�_�_�_ 3_�_�_�_oo&o�_ Jo\ono�o�o�o�o��ׁ  /1_3_\�ATBCKCTL.TM���o+\=;INI9�v5�6%J!0MESSA�GV dqF!�o{ODGE_D� Y&6%�x�O���3PAUS�� !�� ,,		� �� ��4��@�B�T��� x��������ҏ�����B����t�pTSK  �}C?I0�UPDT�pbwd����vXWZD_E�NBbt2*��STApau����XIS$ ?UNT 2�C!�E � 	 �ΝJ�s� �u���yGy�ϻq
�� 
��v5d;C�s��F�А��)�M2��- [\� 8��a��¯��������METr��2i�b# P��AmB`A	4j�@�6w9��@��A�|�٭>a4�>ٸ��>p��5���'>B�>H����SCRDCFoG 1�%1' �^%C"篻��Ϳ߿���<?
Q Z)��e�wωϛϭϿ� &���J���+�=�O�`a���߼1GR��������`NA� ��	4��_ED�`p1���O��%{-�`EDT-�߰�*�B��bE" C���2�
"AO�&
��^����!2��#� �G���� 1��G����6����3��+]���̔(���@Z�l�����4K �������t�&8�\��5�d� ��@���(��6�S0/w��/w/ ��f/���7�// �/C/���/C?�/�/2?��/��8{?���?�f &��?OV?h?�?�?��!9GO�?�O�?i&�pO��O"O4O�OXO��CR ���/__q_ =:_�_�O��O�_"_����NO_�DEL�ߞ�GE_�UNUSE�ߜ�I�GALLOW 1���   (�*SYSTEM�*֣	$SER�V_GR�k_`�pREGhe$�c֬_`�NUM�j�c�mP�MU`֥LA�Y�֬PM�PALap�eCYC10�^�n�`�n%sULSU�o�mr�q�jcL;ttBOX�ORI�eCUR_�ap�mPMCNV6�fap10~�pT4DLIǐZ|i�	*PROGRA�gdPG_MI�n�)�AL�u6� ��)�BT�_n$F�LUI_RESU`w���o��ÄMRvn�`�\�_Β��+� =�O�a�s��������� ͟ߟ���'�9�K� ]�o���������ɯۯ�����#��RLAL_OUT Nk����WD_ABO�Rp/o��ITR_�RTN  �D���ل�NONSTO��Я� 8hCE_�RIA_I,`��������FCFG ���ĨN�o_LIMvb2��� �  � 	��gϳB<�҄��e�@� VϷ��τ�ϨH
��ߒ�2�P}An�GP 1�ޥ�n߀ߒ�>Q�C>  C.���Ef��z���߶Ї��U��Ж�Р�Ъ����Թ������������C���ǀ C�j���J��G?�*�{HE�PONFIπ܎�d�G_P�p1;� �U;ծ�����������,�d�KoPAUS~q1;��� r.�t�;�b� �������������� 0@fL�����6�M��NFO �1?�� �T��B������5Au��9	�]�Ǝ߸@��K �D5Oy����C���($�6�T5+���P� 8�h��Ca��.~�:��1５5��O�ϨG���COLLECT�_�?�x�ǯE�N�p������ND-E�?�;c�R�1234567890'�Bya�/$/&��HC��C)j/�/ y\i/{/�/z[�/�/? �/�/?`?+?=?O?�? s?�?�?�?�?�?�?8O OO'O�OKO]OoO�O��O�O�O_�O�9�ο ��IOG !)�����`�_�_�_�_`WTR6�K2"D](�{Y
�O�^o�#o] jt�i�_MOR9�$;� }��8B���`� �e �i�o�o�o�o�oP�kbb1�:�%pm,t�A?]�]���>q�KFt*�`�R�&�u�tqtrC4  A�j����x�A��*��B�pCd B��d �C  @�r���q�:d�QbZqIJ#'d}?�s9�(pm�����dZqT_DE-FB� {%oR�<�thPNUSE��s����g�KEY_TB�L  ������	�
�� !�"#$%&'()�*+,-./(':�;<=>?@AB�C)�GHIJKL�MNOPQRST�UVWXYZ[\�]^_`abcd�efghijkl�mnopqrst�uvwxyz{|�}~���������������������������������������������������������������������������,����͓���������������������������������耇��������������������4Q��LCKp�ٹ��p��STA���t_AU_TO_DOζkv��IND�ٞ�Rg_T1���T23�pݵʳ��TRL(��LETE��z�_�SCREEN �;�kcsc�*�UʰMMENUw 1)l� <7� @������F��#� I���Y�k�������� ſ׿��6���l�C� UϢ�yϋϱ�������  ���	�V�-�?�eߞ� u߇��߽߫�
����� �R�)�;��_�q�� ����������<�� %�r�I�[��������� ������&��5n EW�{���� �"�X/A� ew����/)\�ʠ_MANUALo�*�DB'a.b�����DBG_ERRL�.�*֫�Q �/�/�/�.L!NU/MLIM���lu�
L!PXWORK 1+֫�/#?5?�G?Y?k?mDBTB_�� ,{-�s�Q�st3QDB_A�WAYT#�QGC;P lr=���"�2�_AL� ٟ�2P"Y�n���lpE(_n  1-�[,p
?POJf�@O}O�6_M�IS�֐�;@�p�CONT�IM���lt��FI
� CMOT�NENDt�DRECORD 13֫� ��OxsG�O�KQ9_x{�2w_�_�_ �_DX�_�_K_ oo_$o 6oHo�_�_~o�_�oo �o�o�o�o�o �oD �ohz���1 �U
��.�@��d� ��������Џ�Q� �u����N�`�r��� 󏨟���;���� &���J�5�C���� ��ȯ7��ׯm�"��� F�X�j��y����Ŀ 3����ϣ���Bϱ� f�տ�ϜϮ���[��� S��w�,�>�P�b�����2TOLEREN�C�4B�B�0L���L CSS_CNSTCY 249%�Y e�B����� �����#�5�G�]�k� }�����������������DEVIC�E 25��  �6o����������������&�O��HN?DGD 6�۬0�Cz9
Q��LS 27Y�8������:��PA?RAM 8,I�2��5&�ySLAV�E 9YE_C�FG :F&d�MC:\��L�%04d.CSV�%@c�B�A &�CH kkO&(/B/X�&2"_!�o/])\!1@JP�Џ#N.A�1n_C�RC_OUT �;Y��1*_NOC�ODz<,G�S�GN ="UR#�M�18-�JUL-23 2�2:00�0A:91�7:51�~� V�hr9n1&�o061�M�����j��1�>��VERSION �):V4.�2.11�KEFLOGIC 1>��/ 	�(1@I��!M�2PROG_�ENB Xa=CUL�S�G `�2_A�CCLIM�F����|CWRSTJNT�G
S���1�MOFLX!2�DINIT ?��"U�ѻ �FOPTu �?	�F�B
 	�R575&'P7�4,Y6-X7-W50QX�4WR2-T�({_�7>
TTO  ]�?t�_�6V�@DEX�G�d�B� �SPAT�H A):A\��_5oGo|�HCP_�CLNTID ?<�6� �+���o��IAG_GR�P 2D� �� 	 D��  D�� D_  B��Т��ff�j�`���o�l��a���%���B�N�C�-�Bz��Bp���e`�imp2�m7 7890123456xq�G�`��  Ao�
Aj{Ad��]AW�A�P��AJ=qA�C33A<�4z1�j�p�!@��]pYA�q��A�����B4�lf�dX�!
�ru�ppQ��Aj�HAeG��A_�pY��AS��pM2�F�RA@(��J���t�J�<�I�@�p��������@��HL��^�p��������33�<��=q@~�R�@xQ�@q��@k�@dz�;@]��Vff؏����� ���s>�l��@e@^J��W
=@Pv�G��@@v�7ڐ.�{d�v���������S�>�M���AR�<(��@5Ґ/\)@_(��@!R�֏  ��$�6��ĭ��� ܯ"�4����V�|�Z� ����<�N������� 0�B�̿R��B�`�r5�༂M�ّe��m>��}R��?�33?9������m7'�����6��4�Fn��L�m@ž�*���ڐ␀N��Z�=@�pAh������c= c<���]>*�H>�V>�3�>�����m<���<�b�a�i�L. ��?� �C�  �<(�UX" 4��>��ё��ٝiA吳 ?�el���t��� �,��H��8�b���r����z����x�?��7��>�(�>!{����=����mo��G��G��m ����I��m����i��@�Ҁ�@Q�?L��Ly�o�g�v\����]p'�@����`8���	�gC� ���Cu��Zl <� ���`�8�O�\���� ��N4\��6{���D5O���K/C��� >T&UP�Q���$��z�	��7E?��;�݈�i ��x�����c��m����6/��dCT_CONF�IG E?i3�eg�%�aST�BF_TTS�G
@UI�#�0�C�A�&� �MAU�@JOJ"MS�W_CFX F�k � �p�:OCVIE�W� G�-�a�� �o=?O?a?s?�?�?�B +?�?�?�?�?OO�? >OPObOtO�O�O'O�O �O�O�O__(_�OL_ ^_p_�_�_�_5_�_�_ �_ oo$o�_HoZolo ~o�o�o�oCo�o�o�o  2�oVhz���@,RC�#{��"!L�~���A�0��e�T����$SBL_�FAULT I��z 8��GPMSK��'��L TDIAG� J\)�!���1�UD1:� 6789012345�p"1�j'�uP&/O�a�s������� ��͟ߟ���'�9��K�]�o�����y��
�>���F&TRECP���
���%���=� :�L�^�p��������� ʿܿ� ��$�6�H��Zρ�������7UM�P_OPTION� ����TR�"�#�����PME�%��Y�_TEMP  ?È�3BȞ 1�s�A.��UNI� ��%1��&YN_BR�K K?6EDITOR����
���_ԠENT 1L��y  ,&�MAI��TLOG� T1��e�&POART2������1��0�&OMAY��[���F��� ��� u���J�����
IRVWAI�����&-BCKE�DT- �/����PICKSIM_ �[���y���$x��� ����������3 WiP�t�������~�MGDI_STAD� !1Ѷy�NC71M�+ C�`�r��
��d�����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S? ��j?|?�?�?�9��? �?�?�?
OO.O@ORO dOvO�O�O�O�O�O�O �O__*_<_�:c?m_ _�_�_�?�_�_�_�_ o!o3oEoWoio{o�o �o�o�o�o�o�o /A[_ew���_ ������+�=� O�a�s���������͏ ߏ���'�9�SA� o��������ɟ۟� ���#�5�G�Y�k�}� ������ůׯ���� �1�K�]�g�y���A� ����ӿ���	��-� ?�Q�c�uχϙϫϽ� ��������)�C�U� _�q߃ߕ߯������� ����%�7�I�[�m� ������������ �!�3�M�W�i�{��� �߱��������� /ASew��� ����+E� Oas������ ��//'/9/K/]/ o/�/�/�/�/�/�/�/ �/?#?=/?Y?k?}? ���?�?�?�?�?O O1OCOUOgOyO�O�O �O�O�O�O�O	__5? G?Q_c_u_�_�?�_�_ �_�_�_oo)o;oMo _oqo�o�o�o�o�o�o �o�_?_I[m �_������ �!�3�E�W�i�{��� ����ÏՏ����� 7A�S�e�w������ ��џ�����+�=� O�a�s���������ͯ ߯���/��K�]� o��������ɿۿ� ���#�5�G�Y�k�}� �ϡϳ���������� '�9�C�U�g�ߓ��� ����������	��-� ?�Q�c�u����� ��������1�;�M� _�q��ߕ��������� ��%7I[m ������� )�3EWi��� ������// //A/S/e/w/�/�/�/ �/�/�/�/?!+?=? O?a?{m?�?�?�?�? �?�?OO'O9OKO]O oO�O�O�O�O�O�O�O �O?_5_G_Y_s?�? �_�_�_�_�_�_�_o o1oCoUogoyo�o�o �o�o�o�o�o_#_- ?Qc}_���� �����)�;�M� _�q���������ˏݏ �i%�7�I�[�u �������ǟٟ��� �!�3�E�W�i�{��� ����ïկ����� /�A�S�m�w������� ��ѿ�����+�=� O�a�sυϗϩϻ��� �������'�9�K�e� [߁ߓߥ߷������� ���#�5�G�Y�k�}� ������������ �1�C���o�y����� ����������	- ?Qcu���� �����);M g�q������ �//%/7/I/[/m/ /�/�/�/�/�/�/ ?!?3?E?_i?{?�? �?�?�?�?�?�?OO /OAOSOeOwO�O�O�O �O�O�O�/__+_=_ W?I_s_�_�_�_�_�_ �_�_oo'o9oKo]o oo�o�o�o�o�o�o�O �o#5O_a_k} �������� �1�C�U�g�y����� ����ӏ�o�o	��-� ?�Yc�u��������� ϟ����)�;�M� _�q���������˯E� ����%�7�Q�[�m� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ���������� /�I�S�e�w߉ߛ߭� ����������+�=� O�a�s������� ������'�A�7�]� o��������������� ��#5GYk}������� �$�ENETMODE� 1NB�_�  �������� RRO�R_PROG �%�
%��an<TABLE  ��L�����<SEV_NUM 
  �� <_AUTO_?ENB  (�9_NO! O�� "  *U�Y �Y �Y �Y � +X r/�/�/2$F�LTR/0&HIS����++_ALMw 1P� ���Y,��+�/2?D? V?h?z?�?�/_�8   �W!�:�� TCP_VER� !�
!Y�?$�EXTLOG_R�EQ�&�))#CSsIZ,ODSTKII�G%� BTOL�  ��Dz�"��A D_BWD��0�@�&�A#�CDI�A QB��C��KSTEP��O�O� �@OP_D�OkO�FACTO�RY_TUN�'d�3YDR_GRP s1R�	�!d 	�?��_{P�*u����RHB ���2 ��� �e9 ����V�{S�_�]{PB����B�CEC���B���A���BFE�]A�]�qA��B���&A���AI��B�>�]�_Wo�Bo{ofo�o�o�o�o � @�:A|=�@9q��o��
? F�5W&b�`��A�ϵ�o	2�o�o\G��]�  v�qA��`�33�r��33�]@UUT��z@�`�pj$>u�.�>*��<�����]E�� F�@ �p&��]J���NJk�I�'PKHu��IP�sF!���]�?�  j��9��<9�8�96C'6<�,5���~����=�����_�� �_&����"tFEATURE SB���@"Ha�ndlingTo�ol 	���E�nglish D�ictionar}y�4D St���ard	��Analog I/O@��I�gle Shi�ft\�uto S�oftware �Update��m�atic Bac�kup���gro�und Edit���Camera�W�F[�CnrRn�dIm���omm�on calib' UI��n͑�Monitor&��tr�Reliaybp��DHCP��]�ata Acq�uis5�^�iag�nos��T�x�oc�ument Vi�eweA�`�ual� Check S�afety!��hanced!�����sʠFrސ�xt�. DIO 1�f�i��&�end��E�rr@�L��B��s�A�rR�1� �@�F�CTN Menu��v\���TP I�n��fac���G�igE��εƐp �Mask Exc���g#�HT��Pr?oxy Svˤ�igh-Spe���Ski�Ŧ�5�m�munic��ons<�ur����s�X����connect� 2s�ncr��sGtru#�qʚ�e���۠J���KARE�L Cmd. L� �ua���Runw-Ti"�Env��^��el +��s���S/W�Lice�nseݣʬX�Bo�ok(Syste�m)�MACRO�s,3�/Offs	ew�V�H5���q�[��MR:�6���Mec_hStop�t��D��V�iS�s���x���T�����odq�wiGtch�ߚӡ�.{��Optm,���'filʬ��gi�V�?ulti-T��Г��PCM fun��Ǣ�o��ޢ����R�egiK�rW���r�iàF����U�Num Sel��� � AdjuG��=�<s�N�tatu��f��Ū�RDM Ro�bot �scov�e)���ea��"�F�req AnlyNW�Rem��5�n7�|����Servo5����SNPX b��x�SN��Clix¡%t�Libr(�DE�� ��W o0�=t��ssag�����0 ��n���0/I|���MILIB�~�P Firm��:�P��Accǐϛ�TPTXm��el�nn����jղo�rquq�imul�a?��bu�Pa�ѱƐZ�(�&�e3v.���ri۠:�USB por[t �iPL�aà~�R EVNT���nexcept����������VC"�rR�I���V��o"��%Wz+S8 SC�4�/SGE�/�%U�I�Web Pl }� >i�'4������x�ZDT App�lP��&?|7Gr{id��playv=(� ���7Rf".7��6����/Y�-10iA�/8L�?Ala�rm Cause�/��ed*�Asc�ii�<�Load�ʠ:JUplP@�l��7�Gu=�rO�BP��Ֆycp�����蠕�RA� �9�gNRTJ�On�e Hel��漿�������1tr;�R�OS Eth
�tڤBeW7iR�$2Dg Pk;�uVIm+�qFd�� �^nsp����Q�64MB D�RAM�O�SFRO��_ېellW��shao gcK�e��Yp�2ltyp�s'��ԗ�B��D�.�ma�iܠ;�T�q�V�R7��FL!PSu�p�c��� pL���cro~���W�4��&���auestz&rtpڡ���/�3DL}�|�Q���Ty,K��l� Bui��n�/A'PLC��uVZ��/sCGl��CRG#�b�$D��@�R�LS[�&�%BUw��%Kі�&�!TA���B�,يE�TCB��ʏ`��/��^�TC���v��%��TEHǟٖ"�ؗV�����/B��F�H����G:� ��n�������H¯���IA߯�ޯ��LN���M��D���D�����N���P��������RR���Sڿ������W.�@Ǣ��$VGFf�x�P2Z���2�H�ǂϔ�B�ϔ�D���Fr�����"TUMT��01J�\�2fߞ\�TBGG��r7ain��UI*ЦU�HMI��r ponU2�8���af{ �R�v>�VKAREL��_#TP� �e��R9� 0�B�o�f�x���� ���������5�,�>� k�b�t����������� ����1(:g^ p�������  -$6cZl� �������)/  /2/_/V/h/�/�/�/ �/�/�/�/�/%??.? [?R?d?�?�?�?�?�? �?�?�?!OO*OWONO `O�O�O�O�O�O�O�O �O__&_S_J_\_�_ �_�_�_�_�_�_�_o o"oOoFoXo�o|o�o �o�o�o�o�o KBT�x��� ������G�>� P�}�t�������׏Ώ �����C�:�L�y� p�������ӟʟܟ	�  ��?�6�H�u�l�~� ����ϯƯد���� ;�2�D�q�h�z����� ˿¿Կ���
�7�.� @�m�d�vψϚ��Ͼ� �������3�*�<�i� `�r߄ߖ��ߺ����� ���/�&�8�e�\�n� ������������� +�"�4�a�X�j�|��� ������������' 0]Tfx��� ����#,Y Pbt����� ��//(/U/L/^/ p/�/�/�/�/�/�/�/ ??$?Q?H?Z?l?~? �?�?�?�?�?�?OO  OMODOVOhOzO�O�O �O�O�O�O_
__I_ @_R_d_v_�_�_�_�_ �_�_oooEo<oNo `oro�o�o�o�o�o�o A8J\n �������� �=�4�F�X�j����� ��͏ď֏����9� 0�B�T�f�������ɟ ��ҟ�����5�,�>� P�b�������ů��ί ����1�(�:�L�^� ����������ʿ���  �-�$�6�H�Zχ�~� �Ͻϴ���������)�  �2�D�V߃�zߌ߹� ����������%��.� @�R��v����� ������!��*�<�N� {�r������������� ��&8Jwn������� � H552���21R78�50J614�ATUP)54�5)6VCAM�CRIdUIFv)28eNRE�52XR63S{CHDOCV�wCSU869)�04EIOC�4�R69XESE�TAWJ7WR6�8MASKP�RXY}7OC�O(3A! (3�`&J6'53�H�(LCHH&OPL�GA0x&MHCR�I&S�'MCS@0�$'554MDSW�!7k'OPk'MPR�l&��(0(PCM|R0g7! 4� �'[51L51�80L�PRS'69`&F{RDdFREQ�MCN93(S�NBA��'SHLEBFM'G�82(�HTC@TMIL��TPA�TPTXYFEL�6� �q8J95��TUTl'95`&U�EV&UECH&U�FRdVCC XO��&VIPdFCSCN�FCSG��IwWEB@HTT@�R6��HCG_WI�GGWIPGS�VRmCdFDGk'H7��R66LR7'Rn�8R53�768�8�2x&R�*4�W66�4R64NVD&R6�'9 �X�9 ֈD0+gF~hCL9IP8KCMS��`n@STY$WTO@�NN`&ORS�&Mv�8OL�hENDuLWS�hFVR��V3D$X{PBV�FAPL�APV�l&CCG@CCRv�&CDWCDL�VwCSB�CSK,6;CT{GCTBHV�p��hC(F�p�xC<WT�C|�ppwTC�wTC&CTE�9�|wcTE�9�0WTF�x�F�hG�xGx�$�H�$�IF��$��GCTUM�hM�M�xN$��P��P�xR�x�hT�S�xW8��VVGF6P�P2 WP2�6e��\�B\�D\�F|V�P��VT��VkTB�wV�IHWG)V�P՗K$WV_V� �)�;�M�_�q����� ����˯ݯ���%� 7�I�[�m�������� ǿٿ����!�3�E� W�i�{ύϟϱ����� ������/�A�S�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ������������ '�9�K�]�o������� ����������#5 GYk}���� ���1CU gy������ �	//-/?/Q/c/u/ �/�/�/�/�/�/�/? ?)?;?M?_?q?�?�? �?�?�?�?�?OO%O 7OIO[OmOO�O�O�O �O�O�O�O_!_3_E_ W_i_{_�_�_�_�_�_ �_�_oo/oAoSoeo wo�o�o�o�o�o�o�o +=Oas� �������� '�9�K�]�o��������ɏۏ�  H55Ȕ��ܻ��R78�50�	�J614	�AT�U�?�5459�6�	�VCAM	�CR�I��UIF9�28n��NRE�52x�wR63�SCH	��DOCV��CSU��8699�0H�E�IOCɛ4(�R6=9x�ESETY�w��J7w�R68�M�ASK	�PRXY���7	�OCOy�3�Y�(���8�3تJ6�7�53(�H�LC�H��OPLGY�0^��MHCR��Sw��MCSX�0��55�H�MDSWٻ�OP�MPR��(��08�PCM��R0`7˅�H���(�51h��51x�0h�PRSvx�69تFRD���FREQ�MCN�	�938�SNBA�ٛ�SHLB	�M�7��ȼ28�HTC�X�TMIL�(�T{PAH�TPTXy�#EL�ʅ�(�8'�%���J95��TUTv�95تUEVx�wUEC��UFR���VCCX�O��VI�P��CSC��CS�GȚ�I	�WEBnX�HTTX�R6ל���CG��IG��I�PGS	�RC��D�G�H7'�R66�h�R7g�Rv�R5�3h�68h�2��R�6�4��66H�R6�4�NVDx�R6�����h�������D0:��FVCLI�g��CMSH�� X�STmY��TOX�NNت�ORS��M��OL��END�Lg�S��FVRH�V3D܈짛PBV��AP�LH�APV�CC�GX�CCRx�CD�g�CDL(�CSBn�CSK�CT��GCTB�� �C8�45 ,C��TC��5 ��TC�TCx�CcTE��� �TE��� ��TF,F�GR,G�-�,H�,IڸE0�,��CTM�M�x,M�N�,PH<P�,R,�TS,W��=(�VGFKP2FX�P2��5@(LB(L�D(LF��VPW;VqT��@(�VTB�-V�IHw�V5��KK��V���_1_C_ U_g_y_�_�_�_�_�_ �_�_	oo-o?oQoco uo�o�o�o�o�o�o�o );M_q� �������� %�7�I�[�m������ ��Ǐُ����!�3� E�W�i�{�������ß ՟�����/�A�S� e�w���������ѯ� ����+�=�O�a�s� ��������Ϳ߿�� �'�9�K�]�oρϓ� �Ϸ����������#� 5�G�Y�k�}ߏߡ߳� ����������1�C� U�g�y�������� ����	��-�?�Q�c� u��������������� );M_q� ������ %7I[m�� �����/!/3/ E/W/i/{/�/�/�/�/ �/�/�/??/?A?S? e?w?�?�?�?�?�?�? �?OO+O=OOOaOsO �O�O�O�O�O�O�O_ _'_9_K_]_o_�_�_ �_�_�_�_�_�_o#o 5oGoYoko}o�o�o�o �o�o�o�o1C Ugy����� ��	��-�?�Q�c��u���������Ϗ���STD�LANG�� � 2�D�V�h�z������� ԟ���
��.�@� R�d�v���������Я �����*�<�N�`� r���������̿޿� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߎߠ���RBT�OPTN���������#�5�8G�Y�k�DPN��� ������������ %�7�I�[�m������ ����������!3 EWi{���� ���/AS ew������ �*�/1/C/U/g/ y/�/�/�/�/�/�/�/ 	??-???Q?c?u?�? �?�?�?�?�?�?OO )O;OMO_OqO�O�O�O �O�O�O�O__%_7_ I_[_m__�_�_�_�_ �_�_�_o!o3oEoWo io{o�o�o�o�o�o�o �o/ASew �������� �+�=�O�a�s����� ����͏ߏ���'� 9�K�]�o��������� ɟ۟����#�5�G� Y�k�}�������ůׯ �����1�C�U�g� y���������ӿ��� 	��-�?�Q�c�uχ� �ϫϽ��������� )�;�M�_�q߃ߕߧ� ����������%�7� I�[�m������� �������!�3�E�W� i�{����������������/ASe��h�������99��$FEA�T_ADD ?	����  	�%7 I[m���� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_o_�_�_�_�_ �_�_�_�_o#o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y������� 	��-�?�Q�c�u��� ������Ϗ���� )�;�M�_�q������� ��˟ݟ���%�7� I�[�m��������ǯ ٯ����!�3�E�W� i�{�������ÿտ� ����/�A�S�e�w� �ϛϭϿ���������DEMO S~   � N�D�V߃�zߌ߹߰� ����������I�@� R��v������� ������E�<�N�{� r��������������� 
A8Jwn� ������ =4Fsj|�� ����//9/0/ B/o/f/x/�/�/�/�/ �/�/�/?5?,?>?k? b?t?�?�?�?�?�?�? �?O1O(O:OgO^OpO �O�O�O�O�O�O�O _ -_$_6_c_Z_l_�_�_ �_�_�_�_�_�_)o o 2o_oVoho�o�o�o�o �o�o�o�o%.[ Rd������ ��!��*�W�N�`� ������Ï��̏��� ��&�S�J�\����� ������ȟ���� "�O�F�X���|����� ��įޯ����K� B�T���x��������� ڿ����G�>�P� }�tφϳϪϼ����� ���C�:�L�y�p� �߯ߦ߸�����	� � �?�6�H�u�l�~�� �����������;� 2�D�q�h�z������� ������
7.@ mdv����� ��3*<i` r������� ///&/8/e/\/n/�/ �/�/�/�/�/�/�/+? "?4?a?X?j?�?�?�? �?�?�?�?�?'OO0O ]OTOfO�O�O�O�O�O �O�O�O#__,_Y_P_ b_�_�_�_�_�_�_�_ �_oo(oUoLo^o�o �o�o�o�o�o�o�o $QHZ�~� ������� � M�D�V���z������� ݏԏ��
��I�@� R��v�������ٟП ����E�<�N�{� r�������կ̯ޯ� ��A�8�J�w�n��� ����ѿȿڿ���� =�4�F�s�j�|ϖϠ� ����������9�0� B�o�f�xߒߜ����� �������5�,�>�k� b�t���������� ���1�(�:�g�^�p� ��������������  -$6cZl�� ������)  2_Vh���� ����%//./[/ R/d/~/�/�/�/�/�/ �/�/!??*?W?N?`? z?�?�?�?�?�?�?�? OO&OSOJO\OvO�O �O�O�O�O�O�O__ "_O_F_X_r_|_�_�_ �_�_�_�_oooKo BoTonoxo�o�o�o�o �o�oG>P jt������ ���C�:�L�f�p� ������ӏʏ܏	� � �?�6�H�b�l����� ��ϟƟ؟����;� 2�D�^�h�������˯ ¯ԯ���
�7�.�@� Z�d�������ǿ��п �����3�*�<�V�`� �τϖ��Ϻ������� �/�&�8�R�\߉߀� �߿߶���������+� "�4�N�X��|��� ����������'��0� J�T���x��������� ������#,FP }t������ �(BLyp �������/ /$/>/H/u/l/~/�/ �/�/�/�/�/?? ? :?D?q?h?z?�?�?�? �?�?�?O
OO6O@O mOdOvO�O�O�O�O�O��O__2]  )XH_Z_l_~_�_�_ �_�_�_�_�_o o2o DoVohozo�o�o�o�o �o�o�o
.@R dv������ ���*�<�N�`�r� ��������̏ޏ��� �&�8�J�\�n����� ����ȟڟ����"� 4�F�X�j�|������� į֯�����0�B� T�f�x���������ҿ �����,�>�P�b� tφϘϪϼ������� ��(�:�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������П� ����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲπ����������0�  1�6�L�^� p߂ߔߦ߸�������  ��$�6�H�Z�l�~� �������������  �2�D�V�h�z����� ����������
. @Rdv���� ���*<N `r������ �//&/8/J/\/n/ �/�/�/�/�/�/�/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?OO 0OBOTOfOxO�O�O�O �O�O�O�O__,_>_ P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o po�o�o�o�o�o�o�o  $6HZl~ ��������  �2�D�V�h�z����� ��ԏ���
��.� @�R�d�v��������� П�����*�<�N� `�r���������̯ޯ ���&�8�J�\�n� ��������ȿڿ��� �"�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ �������  2DVhz�� �����
//./ @/R/d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?�?�?�?�?�?�? �?OO&O8OJO\OnO �O�O�O�O�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�_�_�_oo 0oBoTofoxo�o�o�o �o�o�o�o,> Pbt����� ����(�:�L�^� p���������ʏ܏�  ��$�6�H�Z�l�~� ������Ɵ؟����  �2�D�V�h�z����� ��¯ԯ���
��.� @�R�d�v��������� п�����*�<�N� `�rτϖϨϺ����Ϡ����&�5�:� -�P�b�t߆ߘߪ߼� ��������(�:�L� ^�p��������� �� ��$�6�H�Z�l� ~���������������  2DVhz� ������
 .@Rdv��� ����//*/</ N/`/r/�/�/�/�/�/ �/�/??&?8?J?\? n?�?�?�?�?�?�?�? �?O"O4OFOXOjO|O �O�O�O�O�O�O�O_ _0_B_T_f_x_�_�_ �_�_�_�_�_oo,o >oPoboto�o�o�o�o �o�o�o(:L ^p������ � ��$�6�H�Z�l� ~�������Ə؏��� � �2�D�V�h�z��� ����ԟ���
�� .�@�R�d�v������� ��Я�����*�<� N�`�r���������̿ ޿���&�8�J�\� nπϒϤ϶������� ���"�4�F�X�j�|� �ߠ߲���������� �0�B�T�f�x��� ������������,� >�P�b�t��������� ������(:L ^p������ � $6HZl ~������� / /2/D/V/h/z/�/ �/�/�/�/�/�/
?? .?@?R?d?v?�?�?�? �?�?�?�?OO*O<O NO`OrO�O�O�O�O�O��O�O__&_8Y�$�FEAT_DEM�OIN  =T��hP�=PPTINWDEX][lQ�PP�ILECOMP �T����Q�kRKU�PSET�UP2 U�U��R�  N ��Q�S_AP2BC�K 1V�Y G �)9Xok%�_:o=P�P(oeo;U�_ �o o�oDo�o�ozo �o3E�oi�o�� .�R����� A��N�w����*��� я`������+���O� ޏs������8�͟\� ڟ���'���K�]�� �������F�ۯj��� ���5�įY��f��� ���B�׿�x�Ϝ� 1�C�ҿg����ϝ�,� ��P���t���ߪ�?� ��c�u�ߙ�(߽��� ^��߂��)��M��� q� �~��6���Z��� ���%���I�[���� �����D���h������
3�Y�PP�_ }2�P*.VR:���*�������n PC���FR6:�4�X�T|P|��y�_PI���*#.Fq/��	��<,�`/�STM@k/�/"�/�-O/�/�H�/?�'?�/8�/i?�GIFs?�?��%�?F?X?�?�JPG�?!O�%O�?�?qOF�
JS{O�O��7C��OOO%
Java?Script�O�?�CS�O(_�&_�O �%Cascad�ing Styl�e Sheets�T_��
ARGNA�ME.DT�_��� \�_U_�A�T�_�_}�PDISP*�_���To�_�QNa\o�o
TPEINS�.XML�o�_:\��o]o�QCusto�m Toolba�r�oiPASSW�ORDSo��FR�S:\#�oD`Pa�ssword Configd��� <����+�=� �a������&���J� ߏn������9�ȏ2� o�����"���ɟX�� |��#���G�֟k��� ���0�ůT������� ���C�U��y���� ��>�ӿb�������-� ��Q��Jχ�ϫ�:� ����p�ߔ�)�;��� _��σ��$߹�H��� l�����7���[�m� �ߑ� ����V���z� ����E���i���b� ��.���R������� ��AS��w�* <�`���+� O�s��8� �n/�'/��]/ ��//z/�/F/�/j/ �/?�/5?�/Y?k?�/ �??�?B?T?�?x?O �?OCO�?gO�?�O�O ,O�OPO�O�O�O_�O ?_�O�Ou__�_(_�_ �_^_�_�_o)o�_Mo �_qo�oo�o6o�oZo lo�o%�o[�o ��D�h� ��3��W����� ���@����v���� /�A�Џe�􏉟��*����N��r��������$FILE_DG�BCK 1V������� < �)
S�UMMARY.DyG#�ϜMD:W����ېDiag� Summary�����
CONSLOG��p���ۯ����Console� log���	T�PACCN�v�%�^�����TP A�ccountin�=���FR6:I�PKDMP.ZI	PϿӘ
� ϧ����Exceptio�n$�ջ��MEMCHECK���������/�Memory� Data�����l�)��RIP�E��ϒ�'߶�%��� Packe�t L<���L�$y�e���STAT!���߯� %~C�Status��`�	FTP�������1�mmen�t TBD4�`� �>I)ETHERNEy��f�w�����Ethern�L�3�figura�Cϫ��DCSVRAF(�� �9������ verify �all<���M.=c��DIFF1���)���=�S�diff���t�f���CHG01������C����kv�- 	29 2 ���hz3���K �r�VTRNDIAG.LSw(:�z��� Ope���N� ��nosti�c��.�)VwDEV�DAT������Vis~�Device�+IMG��./@/��/<�k$Imag�w/+UP ES�/�/FRS:\�?\=��Upda�tes List�\?��� FLEXEVEN��/�/�?����1 UIF �EvO�O���,�t�)
PSRBW�LD.CMOϜ�G2#O^?0�PS_R?OBOWELU���:GIG�ϾO�?�O>��GigE�(O~��N�A�)�AHADOW�O�O�O�i_��Shado�w Change������a�)RRCMERRa_F_X_��_���PCFG �Errorq ta�il�_ MA��m�CMSGLIB �_�_�_so�B6e��|0�ico+a�)_`ZD�O�o\o�o��7ZDPad�o l{ )RNOTI���o�ow��Not�ific�� F�AG���՟���� (���L��p������ 5�ʏ܏k� ���$�6� ŏZ��~������C� ؟g������2���V� h��������¯Q�� u�
����@�ϯd�� ����)���M������ ϧ�<�N�ݿr�ϖ� %ϣ���[�����&� ��J���n߀�ߤ�3� ����i��ߍ�"��/� X���|����A��� e������0���T�f� ������=�����s� ��,>��b��� �'�K��� �:�Gp��# ��Y�}/$/� H/�l/~//�/1/�/ U/�/�/�/ ?�/D?V? �/z?	?�?�???�?c? �?
O�?.O�?RO�?_O �OO�O;O�O�OqO_ �O*_<_�O`_�O�_�_ %_�_I_�_m_�_o�_ 8o�_\ono�_�o!o�o �oWo�o{o"�oF �oj�ow�/�S �����B�T�� x������=�ҏa�������,���$FI�LE_FRSPRT  ������A��MDONLY 1�VU�� 
 ��)MD:_V�DAEXTP.Z�ZZ3�䏻�ʛ�6%NO Ba�ck file <���S�6)��� ��@�	�M�v�����)� ��Я_������*��� N�ݯr������7�̿ [�ٿϑ�&ϵ�J�\� 뿀�Ϥ϶�E���i� ��ߟ�4���X���e� ��߲�A�����w�� ��0�B���f��ߊ��~E�VISBCKs�|]���*.VD��|��U�FR:\���ION\DATA�\��w�U�Vision VD� �!�[�m����{�� D�����z���3E ��i���.�R ����A�R w�*��`� �/��O/�s/�/ @/�/8/�/\/�/?�/ '?�/K?]?�/�??�?�4?F?�?;�LUI_�CONFIG �WU����; '$ �3x�{U�=O�OOaOsO�O�O�I%@|x�?�O�O�O__'\ �OJ_\_n_�_�_)_�_ �_�_�_�_o�_4oFo Xojo|o�o%o�o�o�o �o�o�o0BTf x�!����� ��,�>�P�b�t��� �����Ώ������ (�:�L�^�p������ ��ʟܟ���$�6� H�Z�l��������Ư دꯁ�� �2�D�V� h���������¿Կ� }�
��.�@�R�d��� �ϚϬϾ�����y�� �*�<�N�`��τߖ� �ߺ�����u���&� 8�J���[����� ��_������"�4�F� ��j�|���������[� ����0B��f x����W�� ,>�bt� ���S��// (/:/�^/p/�/�/�/ =/�/�/�/ ??$?�/ H?Z?l?~?�?�?9?�? �?�?�?O O�?DOVO hOzO�O�O5O�O�O�O �O
__�O@_R_d_v_ �_�_1_�_�_�_�_o o�_<oNo`oro�o�o�&h�`x�o�c�$�FLUI_DAT�A X���>�a)a�d�RESULT 2�Y�ep ��T�/wiza�rd/guide�d/steps/?Expert�o? Qcu����������Ski�p Gpance� and Fin�ish Setup�D�V�h�z��������ԏ���&h ��`.)`�e!�0 �2`!��c�a6A��ps��� ����ԟ���
�� .�@�R��2oy����� ����ӯ���	��-� ?�Q�)e�)cA�3�E�:W�g�rip*pu� ۿ����#�5�G�Y� k�}Ϗϡ�`������� ����1�C�U�g�y� �ߝ�\�n����ߤ�b��g�%pTimeUS/DST��?�Q� c�u������������
�Enable��(�:�L�^�p���������������� �b�a���������#�24*���� ���1C� �y������ �	//-/?/Q/"�4F\�$qRegionT/�/�/?? +?=?O?a?s?�?�?��America Ͽ�?�?�?OO+O=O�OOaOsO�O�O�)ay�m//�O�/�/#sditor�O7_I_[_m_ _�_�_�_�_�_�_�� Touch P�anel  S (�recommenp)�_>oPoboto�o��o�o�o�o�o�o�L���O�O5�O	_Racces�?���� �����,�>����Connect� to NetworkM��������� ̏ޏ����&�8�J�
�H�^ 9+=S�!_PIntroduct�/���� �*�<�N�`�r����� �Ϻ�̯ޯ���&��8�J�\�n������� ���w�����YVSafet�A$�6�H� Z�l�~ϐϢϴ����� �ϩ�� �2�D�V�h� zߌߞ߰��������� ��ɿ��[�k�}� ������������� �1�C��g�y����� ����������	-D?[(�5��-� �Q����� "4FXj|�M� �����//0/ B/T/f/x/�/�/[m �/�??,?>?P? b?t?�?�?�?�?�?�? ��?O(O:OLO^OpO �O�O�O�O�O�O�O�/ _�/3_�/Z_l_~_�_ �_�_�_�_�_�_o o 2oDoU_hozo�o�o�o �o�o�o�o
.@ �Oa#_�G_��� ����*�<�N�`� r�����Uo��̏ޏ�� ��&�8�J�\�n��� ��Q��uן���� "�4�F�X�j�|����� ��į֯诧���0� B�T�f�x��������� ҿ俣��ǟ)�;��� b�tφϘϪϼ����� ����(�:���^�p� �ߔߦ߸������� � �$�6���?��c�� Oϴ���������� � 2�D�V�h�z���K߰� ��������
.@ Rdv�G��k� ���*<N` r�������� //&/8/J/\/n/�/ �/�/�/�/�/��� �1?�X?j?|?�?�? �?�?�?�?�?OO0O �TOfOxO�O�O�O�O �O�O�O__,_>_�/ ?!?�_E?�_�_�_�_ �_oo(o:oLo^opo �oAO�o�o�o�o�o  $6HZl~� O_a_s_��_�� � 2�D�V�h�z������� ԏ�o�
��.�@� R�d�v���������П ⟡��'��N�`� r���������̯ޯ� ��&�8�I�\�n��� ������ȿڿ���� "�4��U��y�;��� ������������0� B�T�f�xߊ�I����� ��������,�>�P� b�t��Eϧ�i���� ����(�:�L�^�p� ��������������  $6HZl~� ��������� /��Vhz��� ����
//./�� R/d/v/�/�/�/�/�/ �/�/??*?�3 W?�?C�?�?�?�?�? OO&O8OJO\OnO�O ?/�O�O�O�O�O�O_ "_4_F_X_j_|_;?�? _?�_�_�?�_oo0o BoTofoxo�o�o�o�o �o�O�o,>P bt������_ �_�_�_%��_L�^�p� ��������ʏ܏� � �$��oH�Z�l�~��� ����Ɵ؟���� � 2����w�9����� ¯ԯ���
��.�@� R�d�v�5�������п �����*�<�N�`� rτ�C�U�g��ϋ��� ��&�8�J�\�n߀� �ߤ߶��߇������ "�4�F�X�j�|��� ������������� B�T�f�x��������� ������,=�P bt������ �(��I�m /������� / /$/6/H/Z/l/~/= �/�/�/�/�/�/? ? 2?D?V?h?z?9�?] �?��?�?
OO.O@O ROdOvO�O�O�O�O�O �/�O__*_<_N_`_ r_�_�_�_�_�_�?�_ �?o#o�OJo\ono�o �o�o�o�o�o�o�o "�OFXj|�� ��������_ 'ooK�u�7o������ ҏ�����,�>�P� b�t�3������Ο�� ���(�:�L�^�p� /�y�S���ǯ��� � �$�6�H�Z�l�~��� ����ƿ������ � 2�D�V�h�zόϞϰ� �ρ��������ۯ@� R�d�v߈ߚ߬߾��� ������׿<�N�`� r����������� ��&�����	�k�-� �������������� "4FXj)�� �����0 BTfx7�I�[�� ���//,/>/P/ b/t/�/�/�/�/{�/ �/??(?:?L?^?p? �?�?�?�?�?��?� O�6OHOZOlO~O�O �O�O�O�O�O�O_ _ 1OD_V_h_z_�_�_�_ �_�_�_�_
oo�?=o �?ao#O�o�o�o�o�o �o�o*<N` r1_������ ��&�8�J�\�n�-o ��Qo��uow����� "�4�F�X�j�|����� ��ğ������0� B�T�f�x��������� �ᯣ���۟>�P� b�t���������ο� ���՟:�L�^�p� �ϔϦϸ������� � �ѯ���?�i�+��� �ߴ���������� � 2�D�V�h�'ό��� ��������
��.�@� R�d�#�m�Gߑ���}� ����*<N` r����y��� &8J\n� ���u�������/ ��4/F/X/j/|/�/�/ �/�/�/�/�/?�0? B?T?f?x?�?�?�?�? �?�?�?OO��� _O!/�O�O�O�O�O�O �O__(_:_L_^_? �_�_�_�_�_�_�_ o o$o6oHoZolo+O=O OO�osO�o�o�o  2DVhz��� o_���
��.�@� R�d�v���������}o ߏ�o��o*�<�N�`� r���������̟ޟ� ��%�8�J�\�n��� ������ȯگ���� Ϗ1��U��|����� ��Ŀֿ�����0� B�T�f�%��ϜϮ��� ��������,�>�P� b�!���E���i�k��� ����(�:�L�^�p� �����w����� � �$�6�H�Z�l�~��� ����s��������� 2DVhz��� ����
��.@ Rdv����� ��/����3/]/ �/�/�/�/�/�/�/ ??&?8?J?\?�? �?�?�?�?�?�?�?O "O4OFOXO/a/;/�O �Oq/�O�O�O__0_ B_T_f_x_�_�_�_m? �_�_�_oo,o>oPo boto�o�o�oiO{O�O �O�O(:L^p ������� � �_$�6�H�Z�l�~��� ����Ə؏�����o �o�oS�z������� ԟ���
��.�@� R��v���������Я �����*�<�N�`� �1�C���g�̿޿� ��&�8�J�\�nπ� �Ϥ�c���������� "�4�F�X�j�|ߎߠ� ��q��ߕ��߹��0� B�T�f�x������ ��������,�>�P� b�t������������� ����%��I�p �������  $6HZ�~� ������/ / 2/D/V/w/9�/] _/�/�/�/
??.?@? R?d?v?�?�?�?k�? �?�?OO*O<ONO`O rO�O�O�Og/�O�/�O �O�?&_8_J_\_n_�_ �_�_�_�_�_�_�_�? "o4oFoXojo|o�o�o �o�o�o�o�o�O_�O 'Q_x���� �����,�>�P� ot���������Ώ�� ���(�:�L�U /y���eʟܟ� � �$�6�H�Z�l�~��� ��a�Ưد���� � 2�D�V�h�z�����]� o����������.�@� R�d�vψϚϬϾ��� ���ϳ��*�<�N�`� r߄ߖߨߺ������� ���ӿ�G�	�n�� ������������� "�4�F��j�|����� ����������0 BT�%�7�[�� ���,>P bt��W���� �//(/:/L/^/p/ �/�/�/e�/��/� ?$?6?H?Z?l?~?�? �?�?�?�?�?�?? O 2ODOVOhOzO�O�O�O �O�O�O�O�/_�/=_ �/d_v_�_�_�_�_�_ �_�_oo*o<oNoO ro�o�o�o�o�o�o�o &8J	_k-_ �Q_S����� "�4�F�X�j�|����� _oď֏�����0� B�T�f�x�����[�� �󟷏�,�>�P� b�t���������ί� 򯱏�(�:�L�^�p� ��������ʿܿ� ��џ�E��l�~ϐ� �ϴ���������� � 2�D��h�zߌߞ߰� ��������
��.�@� ��I�#�m��YϾ��� ������*�<�N�`� r�����Uߺ������� &8J\n� �Q�c�u����� "4FXj|�� ������//0/ B/T/f/x/�/�/�/�/ �/�/�/���;?� b?t?�?�?�?�?�?�? �?OO(O:O�^OpO �O�O�O�O�O�O�O _ _$_6_H_??+?�_ O?�_�_�_�_�_o o 2oDoVohozo�oKO�o �o�o�o�o
.@ Rdv��Y_�}_ ��_��*�<�N�`� r���������̏ޏ�� ��&�8�J�\�n��� ������ȟڟ쟫� �1��X�j�|����� ��į֯�����0� B��f�x��������� ҿ�����,�>��� _�!���E�Gϼ����� ����(�:�L�^�p� �ߔ�S��������� � �$�6�H�Z�l�~�� Oϱ�s������� � 2�D�V�h�z������� ��������
.@ Rdv����� �������9��` r������� //&/8/��\/n/�/ �/�/�/�/�/�/�/? "?4?�=a?�?M �?�?�?�?�?OO0O BOTOfOxO�OI/�O�O �O�O�O__,_>_P_ b_t_�_E?W?i?{?�_ �?oo(o:oLo^opo �o�o�o�o�o�o�O  $6HZl~� ������_�_�_ /��_V�h�z������� ԏ���
��.��o R�d�v���������П �����*�<��� ���C�����̯ޯ� ��&�8�J�\�n��� ?�����ȿڿ���� "�4�F�X�j�|ώ�M� ��q��ϕ�����0� B�T�f�xߊߜ߮��� ��������,�>�P� b�t��������� �����%���L�^�p� ��������������  $6��Zl~� ������  2��S�w9�;� ����
//./@/ R/d/v/�/G�/�/�/ �/�/??*?<?N?`? r?�?C�?g�?�?�/ OO&O8OJO\OnO�O �O�O�O�O�O�/�O_ "_4_F_X_j_|_�_�_ �_�_�_�?�?�?o-o �?Tofoxo�o�o�o�o �o�o�o,�OP bt������ ���(��_1ooU� �Ao����ʏ܏� � �$�6�H�Z�l�~�= ����Ɵ؟���� � 2�D�V�h�z�9�K�]� o�ѯ����
��.�@� R�d�v���������п ������*�<�N�`� rτϖϨϺ����ϝ� ����#��J�\�n߀� �ߤ߶���������� "��F�X�j�|��� ������������0� ����u�7ߜ����� ������,>P bt3����� �(:L^p �A��e����� / /$/6/H/Z/l/~/�/ �/�/�/�/��/? ? 2?D?V?h?z?�?�?�? �?�?��?�O�@O ROdOvO�O�O�O�O�O �O�O__*_�/N_`_ r_�_�_�_�_�_�_�_ oo&o�?Go	Oko-O /o�o�o�o�o�o�o "4FXj|;_� �������0� B�T�f�x�7o��[o�� Ϗ�����,�>�P� b�t���������Ο� ���(�:�L�^�p� ��������ʯ��ӏ�� ��!��H�Z�l�~��� ����ƿؿ���� � ߟD�V�h�zόϞϰ� ��������
��ۯ%� ��I�s�5��߬߾��� ������*�<�N�`� r�1ϖ��������� ��&�8�J�\�n�-� ?�Q�c��������� "4FXj|�� ������0 BTfx���� �������/��>/P/ b/t/�/�/�/�/�/�/ �/??�:?L?^?p? �?�?�?�?�?�?�? O O$O��/iO+/�O �O�O�O�O�O�O_ _ 2_D_V_h_'?y_�_�_ �_�_�_�_
oo.o@o Rodovo5O�oYO�o}O �o�o*<N` r������o� ��&�8�J�\�n��� ������ȏ�o鏫o� �o4�F�X�j�|����� ��ğ֟������ B�T�f�x��������� ү�����ُ;��� _�!�#�������ο� ���(�:�L�^�p� /��Ϧϸ������� � �$�6�H�Z�l�+��� O����߇������ � 2�D�V�h�z���� �������
��.�@� R�d�v���������}� �ߡ�����<N` r������� ��8J\n� �������/ ����=/g/)�/�/ �/�/�/�/�/??0? B?T?f?%�?�?�?�? �?�?�?OO,O>OPO bO!/3/E/W/�O{/�O �O__(_:_L_^_p_ �_�_�_�_w?�_�_ o o$o6oHoZolo~o�o �o�o�o�O�O�O�O 2DVhz��� ����
��_.�@� R�d�v���������Џ �����o�o�o]� ��������̟ޟ� ��&�8�J�\��m� ������ȯگ���� "�4�F�X�j�)���M� ��q�ֿ�����0� B�T�f�xϊϜϮ��� ѿ������,�>�P� b�t߆ߘߪ߼�{��� ���ÿ(�:�L�^�p� ����������� � ���6�H�Z�l�~��� �������������� /��S���� ����
.@ Rd#������ ��//*/</N/`/ �/C�/�/{�/�/ ??&?8?J?\?n?�? �?�?�?u�?�?�?O "O4OFOXOjO|O�O�O �Oq/�/�/�O	_�/0_ B_T_f_x_�_�_�_�_ �_�_�_o�?,o>oPo boto�o�o�o�o�o�o �o�O_�O1[_ ������� � �$�6�H�Z�o~��� ����Ə؏���� � 2�D�V�'9K�� oԟ���
��.�@� R�d�v�������k�Я �����*�<�N�`� r���������y����� ����&�8�J�\�nπ� �Ϥ϶��������Ͻ� "�4�F�X�j�|ߎߠ� �����������˿ݿ �Q��x������ ��������,�>�P� �a������������� ��(:L^� A�e����  $6HZl~� ������/ / 2/D/V/h/z/�/�/�/ o�/��/�?.?@? R?d?v?�?�?�?�?�? �?�?O�*O<ONO`O rO�O�O�O�O�O�O�O _�/#_�/G_	?_�_ �_�_�_�_�_�_�_o "o4oFoXoO|o�o�o �o�o�o�o�o0 BT_u7_��oo �����,�>�P� b�t�������ioΏ�� ���(�:�L�^�p� ������e��ӟ�� �$�6�H�Z�l�~��� ����Ưد����� � 2�D�V�h�z������� ¿Կ������۟%� O��vψϚϬϾ��� ������*�<�N�� r߄ߖߨߺ������� ��&�8�J�	��-� ?ϡ�c���������� "�4�F�X�j�|����� _���������0 BTfx���m�������$FM�R2_GRP 1�Z�� ��C4  B]��	 ��;�M8E�� F;@ c�5Wo�
�8J��NJk��I'PKHu���IP�sF!�=�{?�  ���89�<9���896C'�6<,5��={A�  /+BH5B�10 !�@�33;"�33¯7]/n-8@UUT�*@9 � {���>u.�>*���<���{>����>��l=<���=�U�=�v�!>1
{:��ܜ:2B8'�Ŭ9IR7�?��9f�͛/$? o/!?Z?E?~?i?�?���_CFG [T �?�? O|O�;NO /
F0HA M@�<�RM_CHKTYP  ��&(�� ROMc@_MsINi@�����@u�T XSSB�3�\� 9�O���C�O�O�5�TP_DEF_O�z��&	WIR�COMh@_�$G�ENOVRD_D�O�F��G]THR֊F ddUdMT_E�NB9_ MPRA�VC]�G�@� �[F@ G���@GAw\H�͊#Iv0�I�ά �?�Oo��o(oK* �QOUUcPAKRK<�@��o�Io�o�o�o��C� � D�o�h1A|A$ B�L.rN�i\�O�PSMTd�Y�*�@t�$HOS�TC�21e�@s���7 MC���T{��� _ 27.02�1�  e�_�q��� ����M�Ə؏���������	anonymous#�Q�c�u�@�������6���� ���F�'�9�K�]� o���������ɯ쟆� 0��#�5�G�Y�k��� ��ҟ���׿���� �1����g�yϋϝ� ���������	��-� p��ϔ����ߺ�ܿ�� �������H�)�;�M� _�q�����Ϲ����� ���D�V�h�z�|�R� �ߑ������������ !3Eh���� �����*�<�N� PA��ew��� �����//<n 3/a/s/�/�/�/�� �/$/?X9?K?]? o?�?��?�?�?�?�/ �?B/#O5OGOYOkO}O �/�/�/�O�?�O,?_ _1_C_�?g_y_�_�_ �_�OT_O�_	oo-o�?o�~�qENT 1�f�y�  P!\�_�o  �p~o �o�o�o�o�o'�o 3\�D�h� ������G�
� k�.���R���v���� ���Џ1��U��N� ��z���r�ӟ������ �ޟ,�Q��u�8��� \�����ᯤ����گ�;���_�"�QUICC0l�H�Z���~�A1�������~�2�����[�!ROU�TER\�8�Jϫ�!?PCJOG�χ��!192.168.0.10��~z�CAMPRT����!��1��#�
��RTu�'�9ߚ� !�Softwar�e Operat�or Panel�w�����`dNAME� !mj!RO�BO���S_CF�G 1emi ��Auto�-started^�DFTP�O�� �O�_���O������� �c_>�P�b�t���� +����������@ \�n��a����x� �����'9 Kn������ ��O�O�O�OV,/� k/}/�/�/�/v�/�/ �/??B/�/U?g?y? �?�?�?�//(/*? O^/?OQOcOuO�OJ? �O�O�O�O�OO�O)_ ;_M___q_�_�?�?�? �_�O�_2Oo%o7oIo [o_o�o�o�o�_�o lo�o!3EW�_ �_�_��o�o�� ���oA�S�e�w��� �.���я����� \n��s������ ��͟ߟ񟴏�'�9� K�]����������ɯ ۯ�0�B�T�f�h�Y� ��}�������ſ��� ����1�T�ֿg�y���ϝϯ�����_ER�R g�����P�DUSIZ  jV�^t����>	�?WRD ?J�7���  guestV�I�[�m��ߑߣ���SCDMNGRP 2hJ�w���7��V�8V�K�� 	�P01.03 8~�   e��?��  ;  �  �� ���������@�-��������x���� 0���y�d����,��>�P�����O  D��d�����������_GROUU��i�������	���5{�QUP��3�������T�YC ����TT�P_AUTH 1�j�� <!i?Pendan��%�`Ϗ�!KAREL:*%.@�KCUewM �VISION SCET����V�K ��J(@:��^p�����C?TRL k�����%V�
4�F�FF9E3�5��FRS:DEFA�ULT3,FA�NUC Web ?Server3*!  5���1�C���/�/�/��/�/?��WR_C�ONFIG l��� 3/��ID�L_CPU_PC�R V�B�8�u0 ;BH[5MINf<!�~y5GNR_IO����V���]0NPT_�SIM_DO�6��;STAL_SC�RN�6 ���IN�TPMODNTOqL�7�;�!RTY�8pu1�6� ��ENB�7���Y4OLNK 1m��E�}O�O�O�O�O�O�OaBMAS�TE�0��aBSLA�VE n��URAMCACHE_��2O��O_CFGI_`CaSUO��l_]R?CMT_OPR �2�ʟSYCLH_{UL _ASG 1o��#�
 �Oo o2o DoVohozo�o�o�o�o��o�o�o�K�RNUMj���
]RIPF_�XWRTRY_CN@�_{U�1���|A���1 ]R�PfRp'^=���=�]0P_MEMBERS 2q���� $�%�r�����w��]0RCA_ACC 2r���  V�4 �E; Z� 3� 6F�s��V�7�S�/P  �`c�U�4�V��5�BUF001 �2s��= �"�u0  u0�1�քJu06x>���Yքvu0F8�.���u0`�qй�u0N�'��u030�B ��ք�ք�Zք�փ�.�.��4u0,I ��Dh�  h����փ��V��փ�Uf�f�(f�7f�UHf�Wf�hf�wf�T��h��f��f��f�U�f��f��f��փ��	��*�9����턷j�y�փ� !׀!0�U&� &�/&�@&�UO&�`&�o&��&�U�&��&��&��&�U�&��&��քք	փ��2��҃ց܁<��r`��� ���������� ����%��-�ց 4�9�=�9�E�9�M�N� T�ց\�a�e�ցl�q� u�q�}�q���q���q� ��q���q���q���� q���q�Őq�͐q�Ր q�ݐq��ց����^����� �2�h�`D�ցL�Q� U�Q�]�Q�e�Q�m�Q� u�Q�}�Q�Q�Q� ��Q�Q¥�᢭����ց��3ɯ҅��� ������­���� ����#���%�3�&� 4�C�B�E�B�M�[�b� ]�k�&�l�{�z�}��� zҍ���zҝ���z�� ��óz�Œӳz�Ւ� z���������� ������&��.� S�6�S�5�S�=�S�E� S�:�U�c�:�e�s�:� u���:Ⅲ��:╢�À:⥢���µ���gQ2�t��4,%&�<ৄ��25�HIS���v�� �S�� 2023-07-18Y&{Ol�~� ��������V)�Y!׀������s!�a�ܚ�U� 9�  ���qY�FXj|� �����1 0BTfx��� ��	�//,/>/ P/b/t/�/�/���/ �/�/??(?:?L?^? p?�/�/�/�?�?�?�?  OO$O6OHOZO�?�? �O�O�O�O�O�O�O_  _2_ �Ƞ/�A�S��_ �_�_�_�_�_�_�����c���d��cO�-�  LU�4�pW iO{Oeowo�o�o�o�o �o�o�oeOPo=O as������ (�'�9�K�]�o� ��������� ���� �#�5�G�Y�k�}��� ��؏�ן����� 1�C�U�g�y����� ��ӯ���	��-�?� Q�?_��T_f_x_���� ҿ����������� ;�;⛳:`񍯟� �ϛϭϿ�������� �+߉�t�a�s߅ߗ� �߻��������:�L� ^�K�]�o����� �����$�6�#�5�G� Y�k�}����������� ���1CUg y��������� 	-?Qcuc��I_CFG 2w�z� H
Cy�cle Time��Busy��Idl��mi�n}�Up|��Read��Dow�� ���Coun}t�	Num �"���`,��7!EQoPROG�xz����p/�/�/�/��/�/?�@USDT�_ISOLC  �z�� O0�J�23_DSP_ENB  B;�c0?INC ys=���P0A   ?� � =���<#��
O1�9:�o ��1�?�?���?O\7OB� Cl3��6"A�G_GROUP �1zB;b<A� �3�	nOO?��/�O��Q�O�O�O�_�O0_B_T_f_���?IG_IN_A�UTO/D�:c0PO�SRE*O<FKANJI_MASK�V��ZKARELMO�N {z�h/��y +_DoVohozo�o�bJ�#|�'~3���e|�_4KCL_L�P�NUMp0�o$KE�YLOGGING��`��bA{5� LA�NGUAGE �z�Jp�DEFAULT Xq6h�LG�}�*��x�0�  }��H  ���+'0�������bƼ���;��
�q(?UT1:\�o� ����0�=�@O�a�x�������(3o��c�LN_DISP ~�?��O�O>��OCTOL9����Dz� K1�1O�GB'OOKq0i}d���������X�|���� ϟ����us�'��	m��yjA%;o��?�1k�_BUFFw 2�B; ���2�����*2ү� � �-�$�6�c�Z�l� ������Ͽƿؿ����)� �2�_π3��DCS ��)�2�1$� c�����������v��IO 2��� 1�3�jA�6�F� X�j�~ߎߠ߲����� ������0�B�V�f� x����������տER_ITM?>d �_?�Q�c�u������� ��������); M_q���I��SEV�`s=�TYP?>.�!3���QRSTt�S�CRN_FL 2��� ��ϧ�����//DTP�p??�C�NGN�AMl4��Jrr�UPMS�GI\�U{5}�!_LOAD'@�G %@*%D�MAYɥ�/G�MA?XUALRM�b�Q�C��{5
�"�!_PR�$�P a�%�� C��i�ٯè�)3H@P 2�w�k �Ʀ	O!t�0��0�P?���2�?�? �?�?���?+OOOO2O DO�OpO�O�O�O�O�O _�O'_
__]_H_�_ l_�_�_�_�_�_�_�_ �_5o oYoDo}o�oro �o�o�o�o�o�o1 UgJ�v�� ���	��-�?�"� c�N���j�|������ ̏����;�&�_�B� T���������ݟ�ҟ����7��'DBGDEF �25?1>1�@�R�_LDXDI�SAm ?+�MEM�O_APg E ?=@+
 d�� ��ү�����,�>��� FRQ_CFG� �27h�A ��@���!�<?4dA%A���R�d�z2�2;��4*z��/�� **:� !���ȟ�!�,�>�k� b�tϡϘϪ���#�25� �����'�� �6�,(��~���lߩߐ��� �������'��K�]� D��h�������*?ISC 1�@)� �)�#��4i�9�$��r�]�������_MS�TR ����S_CD 1������ ��,P;t_ q������ &L7p[� �����/�6/ !/Z/E/~/i/�/�/�/ �/�/�/�/ ??D?/? A?z?e?�?�?�?�?�? �?�?OO@O+OdOOO �OsO�O�O�O�O�O_ �O*__N_9_^_�_o_ �_�_�_�_�_�_o��MKg������&o$MLTARMf���۷Qb ��b��o�dQ�METsPU��b�����NDSP_ADC�OL�ef��nCMNmT�o �eFN�`|�o�gFSTLIw�� ���g~�c��t�ePOSC�F5w�nPRPMl�o�yST�`1���w 4��#�
� ���!��!�#�5� w�Y�k��������ŏ ׏����O�1�C����o��aSING_C�HK  $M7ODAe���Ok�Qn��DEV 	���	MC:�HOSIZE��`ȿ�TASK %���%$123456�789 `�r���T�RIG 1��� lQ�����Lٮ�﯌L�B�YP-�L�Ք���EM_INF �1�ۻ`)�AT&FV0E0���k�)S�E0V�1&A3&B1&�D2&S0&C1�S0=Z�)ATZk�����Hÿ�z�߯Ϣ�A�C���g�Nϋϝ� Q���u��� �����Ͽ@�w�d�v� )Ϛ�U߾��߷��ߧ� ��*������r�}�7� �����������&� �J�\���3�E�W� i�������5�4�� X|�u�e�w� �������0B��f ��EO�{�� //�>/�' �/K�/�//�/�?��/'?L?3?p?�NIwTORPpG ?��   	EX�EC1c�22�83��84�85�8���67*�88�89c�2:" D�2D�2D�2D�2 D�2D�2D BDB�DBC2%H21H2�=H2IH2UH2aH2�mH2yH2�H2�H3�%H31H3�2��R_�GRP_SV 1ݔ@� (w����<� ��>%���6���?�u=���J��_D20�ySION�_DBɐ�͝a�  �p�p�放T =`>�W���PP�PQ�f0N   ��Pf1�X��0�1Qb-u�d1�/oAoSo�aP�L_NAME �!Q�|`�!D�efault P�ersonali�ty (from� FD)�P�bRR�27Q 1�L��XL�x|a�P dzr�o�o�o�o #5GYk}� ��������1�C���2�on����� ����ȏڏ������<]�:�L�^�p����� ����ʟܟ� �[i*��)�:�
)�^�]dP M���������ү��� ��,�>�P�b�t��� ��g�y�ο���� (�:�L�^�pςϔϦ� �����ϫ����$�6� H�Z�l�~ߐߢߴ����������� �2� �F@ G&h� G��]gSP  #�_�q�]bd[�C� ��������D�7�Zj���	���=�@� -�X�N�`�r����������SP�0��	]b-�	`B�<N`:�oA�b����� A�  ��	W�V]`�S �]`��PCT��_s  h���)  �  u$�T&"�C�gy�d���\kR6R �1�ti�P*0 � f2|` � @D�  !?}�#X,?]`<!]aA/��%]d�.]d;�	l,"	� ��pJn �NP`e � � � � �΄ � ��"SPK��K ��K=�*�J���J�?��J9٧�U�p��/SP@_f���"j�@�(E�14!�/�#�N�����;f,1�� �a������-��@¾  T1ÅHZ0Z0� �/�Pc��=��>�]a������l? �?�2-!�3�&.. p�Pm �P���P�  ���P�F�*O�%	'�� � HBI�� �  ����&:�ÈlOß�=��̈́E�"@�O�@�>!�O/K"��&&�&�Q_�  '.T�!-0@2��@����"Z=0@A?C� C�P_C�� Ca0Ce0uCi=%��A�%� 0 �P�l�-hhX�'B�P�Q���A�U]aDz�on?3oo Coio�O�dIA�R�TZ�v�A���  �4@?�ff���o�o�no  #{�!8�@9Gz>L�@�0(!�*(�@uu�0�v�i{!Ht#t$�C?]t�@,���<
6b<߈�;܍�<�ê�<���<�^�Ȭ/�C�A�K"��#,"� ?fff?�@?&&���@�.�8��J<?�\�D�N\��I�R!� -$�)%|�'��
�`$ �oЏ���ߏ��<��'�`�r�]����He�F| ��ҟ����m����J��F�  �F���BG�d GC�qV���R���ů ���ԯ���1��U� @��O���F�IG/�ӿ 1���m��0�B�T�:�9��o�{�33ϩπ��ϸ������{An� ��_�EC��U���<��d�?�؃ߊ�h�߮��I�i4����C CfPa0�¸�Ԑ0؜�@�@I����B>�)A��C�AIA���@�?�\������@ �������=q�A��Ay�I�33@0��@���C�1�������(��Cb��=q��Ů�����H�� G��� G�B�I��(E�� C�e��� I"L�J��HV@G5� E�x C���I3�J0��G���I�� 0 C='�߀�k��� ������������" F1jUg��� ����0B- fQ�u���� �/�,//P/;/t/ _/�/�/�/�/�/�/�/ ??:?%?7?p?[?�? ?�?�?�?�? OO�? 6O!OZOEO~OiO�O�O �O�O�O�O�O __D_ /_h_z_e_�_�_�_�_t�_y�(������r��$e�U���o&o9�3�8�x@oRo9�4Mgulo<~o9ѴVwQ�o�o�4p�+4�] �m�i�o(L:|Ju�P�rP~~�������_�����{R��G�2�W�}�h�  �`��ˏ�� �ڏ����F�4�j�X�p�z��������ԟz����4�"��X�F�|���  2 �F@9�G&h6����9�B�&��L)��C�&�9�@-� �9�o�+�=�O���� ���Ħ�GA�w\]�����ɿ7�?Q��|p9�t�9��9���{�
 ֿ9�K�]�oρϓ� �Ϸ����������#��z����hk�y���$MR_CA�BLE 2�hxO �ћqT�p@����?>𦡆і����кƠ��C���ޱO8�tBǻ���ΝJްޱE�Ҭ޶�ߕ֥�>��š��C�N��|�����a���ް��ER�yx�e����L  ����C֠:�������,bu��(Sѡ"�4��ՠ�y�qBy�ԡ��HE���xlt!�ޱ:�Իv� /ߘ���k������C� �L�>�8�f�\�n��� ����������?��H
�� oq<����ܸ���ܸ�*,** \�OM� �i������޲D�<%% �2345678901i{ f��Rް�ް�ްޱ�
�not? sent 5��WpuTES�TFECSALG&#�egۺ�d.$���
>$���p�޴�޷Y/k/}/�/ �9UD1:\m�aintenances.xml�/��/���DE�FAULTa�\�G�RP 2�M � p��  �%�1st mec�hanical �check�ޱ��z3鰄1�?�� [ph��?�?�?�?�?޲�R3controllerb4,O{?PO���?|O�O�O�O�OAcMY=�O޲"8S!ްQ_��kG8_ J_\_n_�_�JCO�__�_�6/_oo(oh:oLoBC[0geW2�. batter��_�_�_	�_�o�o��o�o_i@dui@ablea50"Pqr�]�g�o������Addg�reas;޷f�B�-ް�#���{@P�b�t�����A
dd�oi�/��+��?��&�8�J�\�AXdj7޶����<ް������
�؟���� �#|too�����>ǟ������ү�A�Overhaul�Ow��"� xް,�3�:5��`�r�������ް$Q�пSV�� O�$�6�H�Z�l� ����߿�Ϲ����� � �2߁�VߥϷ��� �߰�������5ߝ�� k���d�v���� ������1��U�*�<� N�`�r���������� ���&8��\ ����������� �M"q�X�| �����7I /mB/T/f/x/�/� �/�/�/3/??,? >?P?�/t?�/�/�/�? �?�?�?OOe?:O�? �?�?�O�O�O�O�OO �O _OO�OsOH_Z_l_ ~_�_�O�_�__�_9_ o o2oDoVo�_zo�_ �_�o�_�o�o�o
 ko@�o�ov�o�� ���1�Ug<� �`�r��������̏ �-��Q�&�8�J�\� n�������ȟ�� ���"�4���X����� ˟����į֯���I� �m����f�x�����p����5��	 T¿ ���*�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t����޼�  �b�?�w  @�  � ��	�����H�Z�l���*��**  @�>�7����������p,>��e� ^���A���u� ��EWi�Ug y�����/ �/-/?/�/u/�/ �/��/�/�/??��/;?M?_?�/�/����$MR_HI_ST 2�>��0�� 
 \
�$ �23456789C01�?�4�?���?9�)O;O�?$O��O �O�O^OpO�O�O_�O �O_I_[___6_�_ �_l_�_�_�_o�_3o �_Woio o�oDo�o�o zo�o�o�oA�d��0SKCFMAPw  >��0)8�1�`IYu�ONREL  ƚ5rq�0[rEX_CFENB�w
ps�Xu�qFNC��tJOGOVLIM�wqd�3�[rKEY�w���_PANp�x+�'�[rRUN ��,�SFSPDT�YP�x�uZsSIG�N��tT1MOT���q[r_CE_�GRP 1�>�rs�2ڰ9���c�� 8��8&�g����B��� ��x�埜�ڟ�ҟ?� Q��u�,�����b�ϯ ��ȯ���)�;�"�_�������|����7[qQ?Z_EDIT��lw���TCOM_CF/G 1�h}�u��&�8� 
��_AR�C_�r�5�yT_MN_MODE�����yUAP_C�PL]��tNOCH�ECK ?h{ @ ������ ��,�>�P�b�t߆���ߪ߼����ߍ{NO_WAIT_L��l�ՀNT���h{�w��c2�_ERR&߁2�hy�1�6��� ���*��q�����w��O`�g�| E�K��  ��ĜAv��a�Ǝ�@ȴ�i9<O�00 ?���O����p{�Y�PARAuMa�h{�����������1�� = O08Zl Hx���������.��R��?ODRDSP\ã���xOFFSET_�CAR�bψDI�S��S_Aw�A�RK���OPEN_FILE���;���S�OPTION�_IO!�3� M_�PRG %hz%c$*E/W.�WO�[����00��%�d.2  p�v� C�!	 �h�h�!�f���h�RG_DSBL  �7rqK�?eRIENTTO�pe�aC:�prA f�UT_SIM_D�'or��hVlLCT �<�粛$�;��9�ed`7_PEqX���4RAT�� d�u�4�UP� �q>�{ �`OOOBOPI�$���2ރ�L�XLw�x[3�0 C�O�O�O�O�O�O_ _(_:_L_^_p_�_�_��_�_�_�_�_ o�g2 �O/oAoSoeowo�o�o �o�o�oB�o�o 1CUgy�������f�o�~9@�!�N�P�K�]�o��� ������ɏۏ���� #�5�G�Y�(�:����� ��şן�����1� C�U�g�y�����l�~� ӯ���	��-�?�Q� c�u���������Ͽ�s�¯��� �2͠4 A�!S�e�Gυϓ��@�A�����ϭ��� ����!�3�Q�W�u߀����{ ��������	�`����!�x�:�o@1?�Q�c�u��A�  ��V�+��!+�21� 9����s  h��p )  �  u$����� )��&�_�J���^fB�l@O�01���_��� {D��0 ��$  �� @D�  ��?}���X,?+���+�D�����~��  ;�	l���	 ��7pJ3 ������*  � � � ��I � �Ou�H�(��H3k7H�SM5G�22G���GN�3h�`�(ϙ�u�CH50
�R50�����r�û�¾  ��� �� �)��m��AK�µ>+�²���801 io��u����� p m3�P�00� �  � ��u��q�	'�� � "I�� �  �<��o�=���1/C+�@Y/_ Z�!�/��"�����q�9NA0�/  'R0�$t���CA0C����*C. ??�q�pk�Az
b0lw�hhXn�B�� �1��~�p!�5��z n��?3�?�?O.OU/�GD!N2K4a+�����@?�faf�ϏO�O3O �Ј�O�KA8+��OZ>!LS ���J(+�:U��EV^I@99�#?�"T� ,A<
6b�<߈;܍��<�ê<����<�^�q�_�AA�p+���#���?offf?p ?&�P�D@�.�R�J�<?�\�	bN\��U2�Q�@��Ao ��`o�W%�O�o�o�o �o�o�o�o%7" [mD�|�,oNo�Po���xF�  �F��+�G�d GCFQ�T��d��� u�����ҏ������ ��/M��&
��� ���2�������J��O�[�3pޟw�@b�������
<�A3�墚?+�C�����w�)�?��H�O����s�
�4�ț�C���C�࿇�b��xb�a��@I�	�B>�)A�C��AIA��@�?\������ú@� ������=�q+�R!>�I33�@0��@��?C�1���[������C���'��=q�ſ���	H��� G�� G��B�I��(E��� C�^l��I�"L�J�H�V@G5� Eߐx C���I�3�J0�G����I�� E@� C��E�0�i� Tߍߟߊ��߮����� ���/��,�e�P�� t����������� +��O�:�s�^����� ���������� 9 $]oZ�~�� �����5 Y D}h����� ��/
/C/./g/R/ d/�/�/�/�/�/�/	? �/-???*?c?N?�?r?t�?>�(I���^o�pR���5�5����?�?@�3�8�xOO@�4Mgu1O<CO@��VwQ]OoO�4p�+4�] �M�I�O�O�O�O_�LJ:�P�RPC^>�_��l_�?x_�_�_�_�[R�_�_o�_oBo-o  �@�EoWo�o{o �o�o�o_Q��o/{5?uc���?��������A�O�  2 �F@@�G&h6l���@�B���L�ձC��@�@� ��ɏۏ����"�@��oL�^�p�����@ã?���AP@��d�@�@�<���@�
 �����"�4�F� X�j�|�������į֯��?ʶ���-K��y��$PARA�M_MENU ?��E� � DEF�PULSE��	�WAITTMOU�TL�RCV_� �SHELL_�WRK.$CUR�_STYLJ�΋�OPT����PT�B����C��R_DECSNW�4U�� �%�N�I�[�mϖϑ� �ϵ���������&�!��SSREL_ID�  �E]Q�5�U�SE_PROG �%0�%"߇�6�C�CRc�G�]Q8���_HOST !0�#!���ߔ�TTP�߈�ӿ�����4��_�TIMEa�G֯�~!�GDEBUGE��0�6�GINP_FOLMSK]��T�P\���PGA�� |�;���CH���TWYPE-�9�!� �Q�z�u��������� ����
)RM _q������ �*%7Irm �����/��WORD ?	0�
 	PRy���SMAI���R3SUͱ=#TE��S��	��J"COL��Uf)�/��Lc� ��@��`ȯ�dq�T�RACECTL �1��E:� }AP> ?'AP�;P�.�&DT Q屉E0� D � � ��U+0/4	/4
/4/4/2�[QY2�� Y2ԐY2��Y2̐Y2Ȑ*12/4/4/4GЪ12/4/4/2�S �4�5�4�4T���2/2�]4�e4��m4�!�3~3�]4�*e4�m4�u4�F�3)�EF.3�54�=40!T�3N3�U4�]4�e4U�m4�u4�}4�EF��3��4��4��4� �4�p�2Tp�2����2!�4"�4#�4$L/13S�0�3�4��F�3_._@_RY�3��?�5�4�12^3��e4�m4�u4�}4��]4�e4�m4�u4� �V�5�5.?@?R?d?v? �?�?�?�?�_�_�_�_ �_�_�_oo*o<oNo `oro�o�o�o�?�?�? O"O4OFOXOjO|O�O �O�O�O�E��o�o�o �o,t'1Uo��� ������ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� C�U�g�y��������� ӿ���	��-�?�Q� c�uχϙϫϽ����� ����)�;�M�_�q� �ߕߧ߹�������� �%�7�I�[�m��� ������������!� 3�E�W�i�{�����k� ��������%7 I[m���� ���!3EW i{������ �////A/S/e/w/ �/�/�/�/�/�/�/? ?+?=?O?a?s?�?�? �?�?�?�?�?OO'O 9OKO]OoO�O�O�O�O �O�O�O�O_#_5_G_ Y_k_}_�_�_�_�_�_ ���_oo1oCoUogo yo�o�o�o�o�o�o�o 	-?Qcu� �������� )�;�M�_�q������� ��ˏݏ���%�7� I�[�m��������ǟ ٟ����!�3�E�W� i�{�������ïկ� ����/�A�S�e�w� ��������ѿ������#��$PGTR�ACELEN  �"�  ���!��7�_U�P ����2f�n�R�g�7�_CFG �f�SP�!�g�����ĭϸ�I��� � ���{�DEF�SPD ���� �I��7�H_C�ONFIG �\f�N� !�!�5d-��F�  �0�aP����L�!��7��IN~�TRL ɷ�ͦ�8��a�PEv����f�p��,Ѹ�7�LID�����	��LLB �1�� ��M�B<�B4��� M�%��Pպ�� << �?�O�n�O�f���� �������"���<� j�P�r�����8��� ����
Q�@3E�v��GRP 1�����"�@��
����!�AM��D�@ D�@� Cf� @ ��1����	�	,�,��`��uG���´F(BIpP:L��p�!�>�l7>����/.�� =�-=%�T/Q//N/�/r/�/ �/0/�/�/�/?)??�  DzN3W?!�
 >??.?�?�?�?�?�? �?�?!OOEO0OBO{O�fO�O�O�O�J)�A�
V7.10be�ta1�� A���� R�!�A�!��@?!G�Q=wy�#�B���$Q�@����B�l�>4Q@�A���QT �Oi_{_�_�_
FTp���<��_�_ �_�_.� ��O��O� 0oBo,ofoPo�o�A-�p��u0�mf��o@��o���@�AWPl�R�c B��B�>�0uBHfs�d!�2!�PuM���d��)��r�cx�tx�����$|����0��<�-�@�F�0�A�33`��������KNOW_M � �"�����SV ��C�]�m?  ��$��oH�3�E�~��!����M���� �R	��ѐ�lb��^���hhXd��1q� �(�0u8�4�����MR�³��&�oj3�������OADBANgFWD����ST��1 1�f��4�խY�!

��.� _�R�d�v�������� п�'���]�<�N� ��rτ��ϨϺ�����2����	�ݠ�<3���3�/�A�S߂�4p߂ߔߦ��5 ���������6�(�:�L��7i�{����8���������M�A֠��b�O�VLD  ���~�PARNUM  ������죷SCHa� o�
�����	�UPD�����#bb�_CM�P_��d����'��zER_CHK����˒��ƗRSu�ٯ��_M�O֯�_�a�_R�ES_G����
 V_��ch���� ���/
/;/./_/ R/d/7�DT�/ 9oУ/�/�/;���/ ??;�!?@?E?; h�`??�?;���?�?��?;��?�?O;V� 1��vߠ��@�`}\�THR_�INRu�f��d�qFMASS~O Z�GMN}O�CMON�_QUEUE �����
�Qa�N� U�N�F�H SE�NDQ#YEXE._UD BE-P_ SOPTIOW,P�PROGRAM %�J%P<O��~RTASK_Ic��u^OCFG ���O���_
`DATA����kP�
2 ʕyo�o�o�o�olo�o �o	-�oQcu��:oINFO���Wm��DC���� (�:�L�^�p������� ��ʏ܏� ��$�6�hH��w�t�Wl r)l	a��K_a�i�~��ENBd��ҹ�2ԘGa2���� X,		��=��� ���@�N�9�$��8��8�`D��_EDIT� �o����dW�ERFLOXdC�RGADJ �}�A����?
���A�ϦQ�������?�  BzD��ga<8�
�v%$�`\�èr-�g�2����r	H�@lo�cBBP���q@\'�ǽ*۰/ݲ **:�ֿ���q��.@A�� ſ�K�@�c���\I)#Ⱥ��1�[ϩ� g�������w�A.@u� ������O���K�5�/� A߻�e߷ߡߛ߭�'� ��#�����=�� y�s����������� ��k��g�Q�K�]��� ����������C��? )#5�Y��� ���� 1�mgy��� ���_/	/[/E/?/ Q/�/u/�/�/�/�/7? �/3???)?�?M?�?�?�?�?{�	&o0OŠxOWOBD�t$ qO��KEO�OAO�O�O	�P?REF ��Š�Š
ϥIORI�TY�W���ӡMP�DSP�Q��A�7WU�T�V��ΦODUC-T�Q}��O��;OGg�_TG���R���vRHIBIT_�DO���[TOEN�T 1�}� (�!AF_INE�aPog!tc�poGm!ud�6oon!icmX^o�vRXY��}�;�š)� ��o�oŠ��o�e�o :!^EW�{� ������6�H�	*uS���A�J������£>��ѶB�/��z��¤�r��}�A;�,  �P}�8�J�\�n�ť
�߆Zߏ����ҟ��£]�ENHA?NCE �i�}�A�dޏD�+�rV�D�� _SɡӡPO�RT_NUMbS�Š.Uӡ_CA/RTRE���l	��SKSTAaW�[S�LGS`ٸk��;�HPUnothingL�)�;�M��]���������_�T?EMP څY����5q�_a_seiban�OϯO(� N�9�r�]ϖρϺϥ� ���������8�#�\� G߀�kߐ߶ߡ����� ����"��F�1�C�|� g������������ �	�B�-�f�Q���u� ������������, P;`�q����������VOERSI@P�WQ� disab�le^���SAVE� ۅZ	26�70H769'�!4���po�C 		(kR�?;+2/ESeO/x/�/�/�/�*Ag,��/z�n_�PW 1ܸk�20�
B�5<?N?�7�@UR�GE�B�P�^�aWAFz0�QdT�pVW`��4LQ��WRUP_�DELAY �����5R_HOT �%FnQ3�O�5R_NORMAL�8��R
O_O.GSEMI�>OdO�O�AQSKI%P3�p�+3x�O __0_�M�5W_eW O_�_�_�_o_�_�_�_ oo'o�_Ko9ooo�o �oYo�o�o�o�o�o �o5#Ek}�U �������1���U�g�y��5�$R�BTIF�4��RC_VTMOUէå����DCR3��I ��AC��}�C�čC���W?���>��="<��N���`��X	1��$,��H��	��OC�?_ �<
6b<���;܍�>u.��>*��<����U���?����� ��ߟ���'�9��K�]�o��������ER�DIO_TYPE�  !=����ED�PROT_CFG� ��G�4B�H3E���A2�n� ���B� � T�b�����:�����п ��c�ϐO(�G_I�;� Y�[�mϣϑ��ϵ��� ���ߡ���E�3�i� Wߍ�{ߝߟ߱���	� �-�/���?�e�S�� w������������ +���O�=�s�a����� ������������� K9o]����� ����5#E GY�}���� �/�1//U/C/y/�g/�/���/����I�NT 2��9J��ǱG;� ?&;s�x��N?�f�0 l? ~;�/�?�/�?�?�?�? �?OO,ORO@OvOdO �O�O�O�O�O�O�O_ *__N_<_r_`_�_�_ �_�_�_�_�_o&oo Jo8ono\o~o�o�o�o��o�o��EFPOS�1 1�̩  x�/:y�A?c N��x-?y�� ��"��F��C�|� ���;�ď_������ ���B�-�f����%� ��I��������,� ǟP�b����I����� ίi�򯍯����L� �p����/���ʿe� w������6�ѿZ��� ~��{ϴ�O���s��� �� �2������z�e� ��9���]��߁���� ��@���d��߈��5� G���������*��� N���K������C��� g���������J5 n	�-�Q�� ��4�Xj Q���q�� /�/T/�x//�/ 7/�/�/m//�/?? >?�/b?�/�?!?�?�? W?�?{?O�?(O:O�? �?!O�OmO�OAO�OeO��O�O�O$_�Cu2 1��O�O_�_{_ �_�O�_s_�_�_�_2o �_Vo�_zoo�o9oKo ]o�o�o�o�o@�o d�oa�5�Y� }�����`�K� �����C�̏g�ɏ� ��&���J��n�	�� -�g�ȟ��쟇���� 4�ϟ1�j����)��� M�֯q�����ϯ0�� T��x����7���ҿ m�����ϵ�>�ٿ� ��7Ϙσϼ�W���{� ߟ��:���^��ς� ߦ�A�S�eߟ� ��� $��H���l��i�� =���a�������� ���h�S���'���K� ��o���
��.��R ��v#5o�� ���<�9r �1�U�y� ��8/#/\/��// �/?/�/�/u/�/�/"?�/F?,_>T3 1� I_�/???�?�?�?�/ O�?)O�?&O_O�?�O O�OBO�OfOxO�O�O %__I_�Om__�_,_ �_�_b_�_�_o�_3o �_�_�_,o�oxo�oLo �opo�o�o�o/�oS �ow�6HZ� ����=��a�� ^���2���V�ߏz�� ������]�H���� ��@�ɟd�Ɵ����#� ��G��k���*�d� ů��鯄����1�̯ .�g����&���J�ӿ n�����̿-��Q�� u�ϙ�4ϖ���j��� ��߲�;�������4� �߀߹�T���x��� ��7���[������ >�P�b������!��� E���i��f���:��� ^����������� eP�$�H�l ��+�O�s<Y?k44 1�v?  2l��/2/� V/�S/�/'/�/K/�/ o/�/�/�/�/�/R?=? v??�?5?�?Y?�?�? �?O�?<O�?`O�?O OYO�O�O�OyO_�O &_�O#_\_�O�__�_ ?_�_c_u_�_�_"oo Fo�_joo�o)o�o�o _o�o�o�o0�o�o �o)�u�I�m ���,��P��t� ���3�E�W����ݏ ���:�Տ^���[��� /���S�ܟw� ����� ����Z�E�~����=� Ưa�ï���� ���D� ߯h���'�a�¿�� 濁�
ϥ�.�ɿ+�d� ����#Ϭ�G���k�}� ����*��N���r�� ��1ߓ���g��ߋ�� ��8�������1��}� ��Q���u������4� ��X���|������5 1�M�_��� ;A�_��� ��T�x�% ���j�> �b���!/�E/ �i//�/(/:/L/�/ �/�/?�//?�/S?�/ P?�?$?�?H?�?l?�? �?�?�?�?OO:OsOO �O2O�OVO�O�O�O_ �O9_�O]_�O
__V_ �_�_�_v_�_�_#o�_  oYo�_}oo�o<o�o `oro�o�o
C�o g�&��\� �	��-����&� ��r���F�Ϗj�󏎏 ��)�ďM��q���� 0�B�T����ڟ��� 7�ҟ[���X���,��� P�ٯt����������� W�B�{����:�ÿ^� ������ϸ�A�ܿe�  ��$�^ϿϪ���~� ߢ�+���(�a��υ�� ߩ�D��߳���6 1���zߌ���D�/� h�nߌ�'��K���� ��
���.���R����� �K�������k����� ��N��r� 1�Ugy�� 8�\��}� Q�u��"/�� �/|/g/�/;/�/_/ �/�/�/?�/B?�/f? ?�?%?7?I?�?�?�? O�?,O�?PO�?MO�O !O�OEO�OiO�O�O�O �O�OL_7_p__�_/_ �_S_�_�_�_o�_6o �_Zo�_ooSo�o�o �oso�o�o �oV �oz�9�]o ����@��d�� ��#�����Y��}�� ��*�ŏ׏�#���o� ��C�̟g�🋟�&� ��J��n�	���-�?� Q����ׯ���4�ϯ X��U���)���M�ֿ�q�������7 1� �ߧ����q�\ϕϛ� ��T���x���߮�7� ��[�����,�>�x� �����ߘ�!��E��� B�{���:���^��� ������A�,�e� � ��$���H�����~� ��+��O����H ���h��� K�o
�.� Rdv�/�5/� Y/�}//z/�/N/�/ r/�/�/?�/�/�/? y?d?�?8?�?\?�?�? �?O�??O�?cO�?�O "O4OFO�O�O�O_�O )_�OM_�OJ_�__�_ B_�_f_�_�_�_�_�_ Io4omoo�o,o�oPo �o�o�o�o3�oW �oP���p �����S��w� ���6���Z�l�~��� ��=�؏a����� � ����V�ߟz����'�<��8 1�*�ԟ � �����¯ȟ毁� 
����@�ۯd����� #���G�Y�k����� *�ſN��r��oϨ� C���g��ϋ�߯��� ���n�Yߒ�-߶�Q� ��u�����4���X� ��|��)�;�u����� ������B���?�x� ���7���[������ ����>)b���! �E��{�( �L��E�� �e��/�/H/ �l//�/+/�/O/a/ s/�/?�/2?�/V?�/ z??w?�?K?�?o?�? �?O�?�?�?OvOaO �O5O�OYO�O}O�O_ �O<_�O`_�O�__1_ C_}_�_�_o�_&o�_ Jo�_Go�oo�o?o�o co�o�o�o�o�oF1 j�)�M�� ���0��T�:�L�MASK 1�W��N�����x�XN�O  ������M�OTE  ǌ  ���_CFG ���O�l�PL_�RANG ��q[���A�OWER ��W�y�`�SM_D�RYPRG %�W��%����TA�RT �q���U?ME_PRO������H�_EXEC_�ENB  �t\�GSPD��6�>�;K�TDBY�k��RMz�k�IA_O�PTIONQ���^��INGVE[RS��Ȋ
��o�I_AIRPURO� ��Մ1�m�MT_��Tl��`��OBOT_ISO�LCŌ�-�4�0�^o�NAME����n�OB_CATEGňy�փ̀����سORD_NUM� ?q�*��H769  ��t@�R�d�x�PC_TIMEOUTQ�{ xx�S232��1�ȅj� L�TEACH PENDAN���8����Ƽ ��p�Maintena�nce Cons��r����"���t?No Use��� ��@�R�d�v߈�v���GNPOΐ��8�̥���CH_L����^�J�	���!�UD1:1���R��VAIL!�¥��\��SR  ��ʡ8���R_�INTVAL���\��໮��V_D�ATA_GRP �2�ȅ�� D��PL�/�H�S�>� ȅv���n��������� ��������F4j X�|����� �0TBdf x������/ /*/P/>/t/b/�/�/ �/�/�/�/�/??:? (?^?L?�?p?�?�?�? �?�? O�?$OO4O6O HO~OlO�O�O�O�O�O��O�O __D_́�$�SAF_DO_PULS���p[��OSCAN}���[����SCm�����`�Xj�W�p�p
���1�`��վQ�r  H��_oo,o>oPo�_�to�o�o�o�o�o����ib2�d�Qy�d�dq�	�T�i @7�FXjtv&y�: ��t�_ @�sTʠ������T D���+�=�O�a�s��� ������͏ߏ����'�9�K��߯�8w�Z�����n�  =��;�o��ʑ��p����
�t��Di_�jaѰ�?X � ���� �U�Q9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ���������	ߗ���2�D� V�h�zߌߞ߰���� �e�� ��$�6�H�Z�@l�~�����}�0�r ��&�������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�� �/�/�/�/�/�/?? +?������ibk?}?�? �?�?�?�?�?�?OO 1O?IROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_��_�_oo&o8o,x� a��Co�o�o�o�o�o �o�o�o"4FX j|���zmo�\��v��+�����	12345�678]2h!B!��%�\1}�k`�T�f�x��� ������ҏ��lo� �1�C�U�g�y����� ����ӟ���	��-� >���a�s��������� ͯ߯���'�9�K� ]�o���@�R���ɿۿ ����#�5�G�Y�k� }Ϗϡϳ����ϖ��� ��1�C�U�g�yߋ� �߯���������	�� -���Q�c�u���� ����������)�;� M�_�q���B������ ����%7I[ m������� �!3EWi{ �������/ ///�S/e/w/�/�/ �/�/�/�/�/??+?@=?O?a?s?�?McE��?�?I/�?�?O�Cz  BpIj_   �H2_b� } �6F
[G�  	�AD�?�O�O�O�O�KDo�<�uO_$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Voho�O�o�o�o�o�o �o�o
.@Rd v�������D#��B�1iA�<�� �iA  �/�I��v,�mA>mAt  6@m�����x`�$SCR�_GRP 1���*P�30� �� ��A ��	 Ё�؂�� �1����w��#��J��M�K@G�DC�v���N�G��L�	M-10iA/�8L 12345_67890k@��� 8k@MT20� ͐-C
ș�X��A^H �؁�Z�ǁ'�ǁ�C�G���-�	�v����������ά��H�؀_�܇ǂ���@�5�G���o�A"����������^� �h@,V�- � �B�%@Ɛ������A6@ � � @�@8��N�?��^���H%@q�K��F?@ F�`�£� ���ϲ�������!�� E�0�i����8�h�0ߑߣߵ�B���X� 	���-��Q�<�N�� r���������O� q�3�!�F��]@C��x��B`�8�>����~�6�i�@8���%@���ȗ�'��?�-DA��1a�]�$> �A2�A T{��
i���� (� �  $��H3l)J��Γ���ECLVL  ��A��7�?A���*SYSTE�M*�@V9.10�214 �8/2�1/20�A ��@�z�SER�VENT_T �  $ $S_�NAME !^	 PORT�@!�ROTO! �_�SPD  ���/ TRQ  � 
,#AXISr5!:'2  2c��,#DETAIL_�  l $?DATETI! ERR_COD�#IMP_VEL4@w 	�"TOQ�$�ANGLES�$D�IS��&" G%%o$LIN�" ,#wREC5! ,!tO%i � MRA�!� 2 d2I�DX!��$B  ��0$OVER_LIMI I ـ�,#OCCUR5!�  �+COU�NTER�"+ FZ�N_CFG5! �4 $ENAB�L�#ST� "FL{AG"DEBU�3�R�!�~3��5! �� 
$MIN_�OVRD�@$I��� �2�1�5FAC�Ee"�1SAF�7MIXEDL�9�!�2�ROB%$NE�&APP�"�SHE�LL�4	 w5$J?@BAS�#�RSR_�5  ?$NUM_y@� � xA1�'y@2��J3�J4�J5�J6ʜJ7�J8�'lARO�O � CO�ON�LY�$USE�_AB#xBAC�KENB�  PIN�>0T_CHKSO?P_SEL_�0,Yg_PU;Qo1M_�!;OU#PNS|F P�YC�&�0EPM�%TPFWD_KAR�!� P�!RE$$O�PTION�2$QSUE�Y" D�RYRB�$CSTOPI_3AL;SYCEX+STQl�P�$XTSPM1i�2"MA�1STY�;TSO
`NBRDIGQTRI�3�Q�W�INI�M& 8bNsRQxf`ENDNd�$KEYSWI�TCH�S�QZa�TH}E�PBEATM�SPERM_LE�"R�QE� �gU�SFd��RS_dDO_HO�M�0ORA/PEFP0 !"0�3U ST�bR�C�`OM�#�!OV�_MSJQ ET_IOCMN+S�W5a���XEHK !
 gD �7qSU�"f�RMP+S� PO7B�$FORC�SW�ARNQ�2ZCOM�rP 7�$F'UNC��3U	0}QSAR'`�u2�v3�vQ4�q�2C0O�PL�ry�"�XUNLOeP��$:�ED� ���SNPX_AS�2 0�@ADD|�0�1$SIZ�!�$VAR�'MU/LTIPRZ��p�A�q � 1$tY[�r	�B`��"�AC� ΆFRI	F">0S�P�y"t���NF{dODBUS_ADw2�B��&�CM�aDIA�q$DUMMY15ajM�3J�4J��Sz@>  � x��"�TEqM�8J�SG�L��TAJp  &�0���@J������STMT�Q��PS3EGb��BW�P���SHOW��!BA=N̐TPOF�M��9J�0J�(a+ V�C�G�2 ��$�PCpP?0-�G3$F�B�qPD�SP�PA�FPF�L VD/��2�� ��!A0 ��@� ���p���p��P	������5��6��U7��8��9��A��B���p��h ��Ր��F���P���T�P����l�P�̩1٩1�1��1 �1�1�1*'�14�1A�1N��T!ǘ�2��2��2��U2̩2٩2�2�U2 �2�2�2'�U24�2A�2N�3��U3��3��3��3��U3̩3٩3�3�U3 �3�3�3'�U34�3A�3N�4��U4��4��4��4��U4̩4٩4�4�U4 �4�4�4'�U44�4A�4N�5��U5��5��5��5��U5̩5٩5�5�U5 �5�5�5'�U54�5A�5N�6��U6��6��6��6��U6̩6٩6�6�U6 �6�6�6'�U64�6A�6N�7��U7��7��7��7��U7̩7٩7��7�U7 �7�7�7'��74�7A�7N��V�P�`U3" �< �B
)�� !� x $TOR��Q@�  �"M$ RX1 L@BQ_W0R�P�%T!�p�$S[C�Q�p�_U�����*0YSL�   � x���7���m��0���`�R�VA�LU�5QP�V]�F��ID_L�"%H�I*I�r$FILcE_xSM$BD$s�}0�SA21 �h5y E_BLC�K�S�"���(D_CPU�)y��)m��3P/�b$p"�`sRR ? � PWY0Pl�� 1LAƑS11�314RUN_FLG(54,14�`/5M14M15HrP4o0�4W�T2�Q_LI��r  k@G�_Ob�PP_E3DI+R��T2 @�3�20�$P�!�����TBC2x� �}�8P/0T�Q�1�FT'dD5cTDC"/0A`a�0@M	�FL.AGTH���DD�OPGRQH��pERVE(crD5crDa��0�BC4PG@ �X -$�ALEN`(c�D5c�@`RA�PLF��W_k�#1�A�:$2�GMO�!C�S�DPIZP�F!Y8̝@![DE1U�LA3CEXrfCCB���`_MA^�0VjU@W�jQTCVq\�Q@WT �a�Z�U�Zd�/S]��UT@S]�J@`AG�M�T" Jjgv�/Ua@U�A2)pp\�5a.S6H�JKHfVK$�ZaU�Zaa�O`J�ra^c�JJfcJJncAAL^c�`fc�`�fm��b5OC�PN1�\�`�[nP�L
P_�� oqv�0CFb� `5GROU ���P��N�0C�� pREQ�UIR]B�EBU�̓�A�V$T1P2�Vq�@@v�1a��4� \�p�8APPR�LpCL�
$�0NN�xCLO�0�yS:E�y/U
�1�� ��0M,@oP�PF��t_MGI��pCx�z ��d�lP�BRK�N�OLD��RTM!O�1I�6��uJ�0H�P�dLPfcLPncLP�c(LP�cLP6��7�������A�4�# Ir�B$��U��PATH���� ��H��p[p�.��SCA�2L��r�qI�N�BUCP�A\�C�f�UMe�Y�@�  `l�&!xA��������~��PAYLOAD��J2LR_AN$AȓL0ҙΑޑ��R_F2LSHRlD�LOӔ[���i��i�ACRL_@�AY�L�U���gbH�΄$H�z�FL�EX�s�1J�6 P�r�?
OqO�Om"|���E  :�O �F@P�#��Oha@P�O�O�LF1#�q����O@__0_B_T_��E^_ p_�_�_�_�_�_�_�_ �ȩ��WcHd����o�!o3o"�:jT�Ǌ�X raFe���QeZ�3� ]ooo�o�`�e�e�e�e��o�o�o�i�BJt! ��0#5 cAT��Hq�PEL��T1p�OxJ[p VpJ�E3�CTRU���T�N)l�@wHAND_VB��� ׄ7" $��F2�<D��SW�g�v#� $$M��yM #��2�-�O� �q�K��A) ���v(!h� �A(��#�A1�A@�s��� #�D1�D@�P2 �G"0		ST%�42�NC�DY.0�p �T�{����@�#������Hg��K�-�G�P ��������������ʂs 	��ׄ$ ���� Ʊ�qOASYM0��IpB0�#wL��P�_n0 A�a�t�^�`��~�������ƓJ͜~�ߚ�������_VI��x<(�sM V_UN�2; b#��
�JIez"� z"�~$4��$�&=��P@P�~�_�q�5;������ς�0HR�0�1a%��01���2DI@��;sOO4��10�&) �Ђ�IeA��4��|1����3��|�����20 ' � -��ME���Х24�"�TC0PT����1�`�d����8��1�9T��a $DUMMY1���$PS_��RF�^�  �(F�pFLApYP2�BB�3$GLB_T� E5]E�0��р۰��1�( X�p@wׁST���VpSBR�M�21_VRrT$S/V_ER�O��C��CCLw@�BA�Ol2,0GLD EWq�) 4p�1$Y
��Z��WS>`���A�0e���AU�E*� ��N P�$�GI��}$�A �)�CPq+� LpAV�}$Fz�EIVNEAR��N��F�Y�TAN�C��2 �JO�GR�t� ,�?$JOINT=�Nм���AMSETq-�  >WEvU�:�S�A��p]R;�q.�k ��U��?�VpLOCK_FO����K0BGLV��G�L:hTEST_X9M�p�QEMP�PRrq^buB%`$U젌�B=�2*VpS�a+�Ob��*`�a)�ACE��`RS�` $KAR�P�MQ3TPDRA8�@�d�QVEC4��fֽPIU�a,�aHE�,`TOOLe��cVvd�RE�`IS3�rr6����ACH�P�[p-qO>��3D3ړ�QPSI�r � @$RAIL_�BOXE=��@R�OBOUd?��AHOWWAR��tq%@@qROLM0B�u ��=t�r0�bp��ـO_�F1�!�@HTML5D1U�0@�B2q�ځ/�_	�R�`OB��0�r]��Q�p�F;OU�R1 d�@�e�)�v�P�%`$PIPVfN0�rbr2q𫰄a�p�CORD�ED*`6���PXT$V�DQ),0,�O�0�Q7D \@OB��z� *`����C[@���|�wSYS��ADR{��,0�0TCH:� 73 ,��EN52��A1a_AT�	�{nd,0VWVA�1?4 � �`�B�E5PREV_RT~�$EDITT�_VSHWR1��F(s�� Q< D�0������$HEA�D�� ���\�K�E Q@CPSPD.��JMP��LD5��R�g45������I_`S{�C��NExp|��TICKe��oM���1�HN�A6 @����Ñ_GPR�Yv��S�TY	�>qLOwA���N� �7 t 
�O�G�%$4�AT=:�@Sq�!$p!=А�1HEy0GFPRR�S�QU�`X�IB;!TEsRC�03��TS�8 HP�@.�0�-���a^�O�0�3���IZJDAQFE$AP�R��1Ap���.�PU�Aဵ_DO�R�XuS�PKD6AXI���s�aURI��|� {p@�͆��J�_�`߂�ET�P3b��5���F5��AB8�D9Hw��!@�S=R��9l �� M�%�[�8�m�K�[�V� [�d�[�t��Ŗ��Ŧ� �Ŷ�����������!��C6���C�ͯ����YQSSC_@ o: h�@DS`���a@SPv0��AT���L���?��BA_DDRESsB_��SHIFA�{`_2+CH{�ɁI~@���TU~@I*� };�rCUSTO�*aVbIj2< �Gh���d�
^j
�rV8-����0= \�@G�A���o�>��P��C���A��~�F��B���T�XSCREE��>z<0��TINA�COP��AT�A���? T���@d�߁�A��@L���ނ��H�[�RRO �Pހ��E�4v��UE�@ �-���6@S�A߁RSM?���U��
�D6��00S_S��i�������i�Cb��3� [2?��UEAp2��Bp�GMT� LҜ!���@O�U �/BBL_BpW�0�0�B ���vOQ�LE�zpE��RIGH�BRD<�D�CKGR�0��T����WIDT�HHs���2!ABAqo�UI�pEY�Ђ�1C6��p�p��bpl�BACK��0B1��A�0FO�DL[AB��?(�0I@p#b$UR�qq-��
�0Hl� D 	81�P_����0R P%b/�Hx A���)O�0EI��G� �U� �R3b�qLUqM�Ķ�ERVM���@
P�PF�0�GEu{Q�������LP4%
�E���)�Q'��_(��_(,p^)5*\+6\+7\+8A"�@�3k��P��F,qa�S�PE	USR��DG <�@�0U�ERT�ERFOB�ERP�RI�mLp�!30T�RIP^qm�UWNDOg5H<Pà L0���q��|aްؠ� I�� o�G ���T�p�� �2O	S�1�6R�r�v3�a�AJ�OS^�2b��p{bU<!�AK�?�?��8<"a�v3OFFT`�@�L�@�3OU@ �1J�@?DgDK�@GUفPfA��C}ьG�SUBb��@/ SRT�0B�MI��Q�p�O�ORBp�ERAUDT��DT�I��A_R���N |]��OW�Ny0�$SRC�}�����DT`>UR�M�PFIy�y��ESP|�G��u#��'�ru1Rm�6O `&@WO���=��7COP!A$հ{0�_YPr�Q.��UWA_�Cra�Q�P�S�Qrp��4��rW� P?�?SHADOW��s~"a_UNSCA�c8"c�/cDGD7q���EGAC�Sd�O�P�PG�Q���STE���O��t�kPE"��VWDt�TRG�6R� �>��jMOVE8}����bANG���f�-C�f�3�bLIM_X!Cv'Cv�hq|���g?06��`��VF8���C}VCC���5S?�C��RA���`�ϥD��@NFA�R�@�]�E,�Q>0G�����R:�{0DE�c�p���p6T�# i�؁ϣ�u��㡹W C% �DRI�`��aV[�*���S�D�$MY_UBY�$�}�3ϥ~���b����a��P_8`�y���L��BM��$�DEY
�EXXc ���UMUِX�d�����US��˰.0_AR�"B#06��fG�PACIqt�`HQ�d�I�-CI��3I����QR!E���1f�sI�N�U ?�PG�`!P�⎐G0�sR�0�AV�k���B	�R��R�dSWA�osh I��n�O�!�A��[�E� U���ah Yt0�sHK��W����aS���Q��cEANS��P���0�r�MRCV6X ��- O�pM�C��	p��?C����REFb ������
r�ِ0���ꡨ�꡹����A�_ ;PW�B�o����`��k��\���r�A�r3Y ���a��ϒ�1`�$GROU���3��H¶�s�pT����20a$ ����0X V�Ӱ��ֱ���UL�qW2�PC%p�X��NT�S+�b*��6��!6���L��_Ű�_�(�k��!�pTIЙ��Z t@MD�@A�P_HU�q�`��S]A�cCMP}�F��(���Ų�_��Rqty����W�j�X�ɗQVG�F`S[� ��M0����UF_`{�˂��@JʼRO� �T�շ����|.�UcRE9��6�RI;���I&༨�o�o{FQ�yFQ'C`wIN�H��xx� V�1,r��A��?�W�|��Q/��V큂��LOp'�\apx �����!NSI"�VIA_�R;�\ }�� HDR )�$JO� b?�$Z_UP)p��Z_LOW������ �\(p���P鱬3 �9���Ⴐ��'Q�����"�]� 0��PA� �CACH���}����P��!�P]SC(qIBӉF#���T� ��|�$HO�1R��/�%� "f������?�RQ0!���cPVP��� H_'SIZ�sRZ��M0��N�Q�MPr
�q�IMG�d��AD�	�RMRE���W7GPM�pNDRP�VASYNBUF�VVRTD� W��?OLE_2D,t�c�1@C�qUۃ��Q���ECCU{�V�EMe�}�d��VIRC��
" {��LA��RQ}0\0��AuGR�XYZ)��C�W�������A2�T�p܂IM���G`��GRABBB�1Y�b�p ���^�p}
�CKLAS�p�b�Y@_  񱒵�T��5P@�21T$8b��p!�` ���SP�G�%TQ�RQ�q�P��"x�I�$|��=�B?G_LEVE�QL��PKL��"ѥ�GI�� NO�Q܁+�͐H�ObPRa �  �F����E6S��g�]2RO�cACCE0e@����x4VR�A`�y1܂R`� AR�c�PA@�>��D�SR�EM_BQ$'0�"J�MPU�XAbi$1�$SSlSFD�Ќ"��|�Y@c  ���S� ��N/D,�LEX�&dbSdqg`��&DR�w$YQqH(`hqH҄�c��P2h��e� �є`V|��cPMV_PI���DX�`�@3����IF&�\rZ�JT�E�@��0�H���E�AGAU?��LOO�d?�JCB�TZ�'B`H +cPLCAN'r��L2��Fw ��D?V5Y �WM��~Ppu�T�FS��U�Q �ѥU����V2DbX9�1LRKEZq�1�VANC]C ��VR_O�|`f (�p8�s$\�3Zr��R_A3� g 4��dovn#p� �B��h h��9��\ĬvOFF�sfW@X�����EA��
� LSK��MN��q�g S`��|@c"i� < WJ��=�UWMMYY���\��D�P�	@CU���1�U�pj $��TITV1$3PR8A��OP����SSF���Cki �|t6���`�SMO!�l%BXC�4J�p��;ZD�vm DQx�AL^1IM; ��0�IN�MSG_QB�Sw7 �_��pn%B�w��%�M�� �XVR"�o�I"�pT�5$�Z7ABC��p��Ƃ���Ӡ
�@%��`V�S.� q � �w0��=�CTIVeAIO�b�	�s�ITVLW�DV�@
l�"��2� DI�� @����|A��d�p��N�LSTs�p��ݰ��_ST���(1%�DCSCH��r LQp������~P1��m�W GN�����r���_FUqN�� �1ZIP!�Ss%B� L8�L|��ѢAZMPCF�ʅt�r9���L�DMY_LN$pq���M&�˄u �$��Q�CMCM���CLCART_���P�a $J����D=��¢ ��u�ǥu���_�p����UX�P�UXEUL����
��̥
��.��>���FTF���k������v �*� �Q`��Y%�D.  w 8 $R� yU�Q��EIGHe3F�x?(�0��0��`��A$x �=0�sqF�$B�����b�_SHIFB�	�ReV�PF��1�	$)��0C�ঢ���d�pl� �r�"l��D|ȕ��C �NV�a���SsPH�0%�y ,�0���ֿ��$S{0D�EFAUn�B���?������'HOT�������MIPOWERFoL  �� �Ž%�WFDO��� �� ��Y��`1 ����q�� �L!ip_EIP�5ԑ����j!A�F���`�߼�!F�T�������!���-����S�!ER9MHQp�7�B� ��f�@o�5黎���!OPCUA������7�!T!PP�@8���d&����!
PM�p�pXY����er���J�����f��!RDM�-@V��g
g!OR90h��hV��!
h�~�����i���!RLSY3NC &8�K�!ROS��r�y4:�!
CEL�#MT�`���k���!	��PS���l��//!�WAS�RC6��m/{/!��USB|/��n|j/�/!STMP��/��o�/?�7?*�?`=e�I��KL �?%q� (%SVCPRG1`?D�:�52�?�?�03�?D�?�04�?�?�05 OD%O�06HOMO�07pODuO�08�O�O�09�O�K�4~�O�1�?_ �1�?=_�1�?e_�1O �_�1:O�_�1bO�_�1 �Oo�1�O-o�1�OUo �1_}o�1+_�o�1S_ �o�1{_�o�1�_�1 �_E�1�_m�1o� �1Co��1ko��1�o e?w2�0~?�00�u��1 y����������Џ	� �-�?�*�c�N���r� ����ϟ�����)� �M�8�q�\������� ˯���گ���7�"� I�m�X���|�����ٿ Ŀ�����3��W�B� {�fϟϊϱ��������k:_DEV ~q��MC:��4���GRP� 2q����0b�x 	� 
 ,c��|�<�hߥ� ���߰�������#�
� G�Y�@�}�d���� ������d�1���U� g�N���r��������� ��	��?&cJ �������� �;M4qX� �����/�%/ /I/0/B//��/�/ �/�/�/�/�/�/3?? W?>?{?�?t?�?�?�? �?�?O�?/OAO�/eO O�O�O�O�O�O�O�O �O_ _=_$_6_s_Z_ �_~_�_�_�_�_HO�_ 'o�_Ko2ooo�oho�o �o�o�o�o�o�o#5 Y@}dv�
o �����1��*� g�N���r�������� ̏	���?�&�c�u� ���P���ϟ���ڟ �)��M�4�q�X�j� ����˯�����%� |��[���f����� ��ٿ�������3�� W�i�Pύ�tϱϘϪ�\��7�d ���	�� �	�B�-�f�Qߊߙ��%��߾�>�����у���������� �9�'�]�k�ߐ��� S������������ ;�}�b���+������� ��������C�i�:y� m[����  ?�3�Ci W�{���� /�///?/e/S/�/ ��/�y/�/�/?�/ +??;?a?�/�?�/Q? �?�?�?�?O�?'Oi? NO`OO9OO�O�O�O �O�O�OAO&_eO�OY_ G_i_k_}_�_�_�__ �_=_�_1ooUoCoeo goyo�o�_�oo�o	 �o-Q?a�o�o ��o�����)� �M��t��=���9� ��ݏˏ��%�g�L� ����m�������ٟ ǟ��?�$�c��W�E� {�i�������կ��� ;�ů/��S�A�w�e� ��ݯ¿Կ�������� +��O�=�sϵ���ٿ c��ϻ�������'�� Kߍ�r߱�;ߥߓ��� ��������#�e�J�� �}�k�������� +�Q�"�a���U�C�y� g����������'��� ��+Q?uc� �������� 'M;q���a ����//#/I/ �p/�9/�/�/�/�/ �/�/?Q/6?H?�/!? �/i?�?�?�?�?�?)? OM?�?AO/OQOSOeO �O�O�OO�O%O�O_ _=_+_M_O_a_�_�O �_�O�_�_�_oo9o 'oIo�_�_�o�_oo�o �o�o�o�o5wo\ �o%�!���� ��O4�s�g�U� ��y��������'�� K�Տ?�-�c�Q���u� �������#����� ;�)�_�M���ş���� s���o�ݯ��7�%� [�������K�����ſ ǿٿ���3�u�Zϙ� #ύ�{ϱϟ������� �M�2�q���e�S߉� w߭ߛ߽��9�
�I� ��=�+�a�O��s�� ����������9� '�]�K��������q� ��������5#Y �����I���� ��1sX�! �y�����9 /0/�	/�Q/�/u/ �/�/�//�/5/�/)? ?9?;?M?�?q?�?�/ �??�?O�?%OO5O 7OIOO�?�O�?oO�O �O�O�O!__1_�O�O ~_�OW_�_�_�_�_�_ �_o__Do�_owo	o �o�o�o�o�o�o7o [o�oO=sa�� ���3�'�� K�9�o�]�����̏ ������#��G�5� k�������[�}�W�ş �����C���j��� 3�������������� �]�B����u�c��� ���������5��Y� �M�;�q�_ϕσϥ� ��!���1���%��I� 7�m�[ߑ��ϸ��ρ� ��}���!��E�3�i� �ߐ���Y�������� ����A���h���1� �������������� [�@�	sa�� ���!�� �9o]���� ��/�!/#/5/ k/Y/�/��/�/�/ �/?�/??1?g?�/ �?�/W?�?�?�?�?	O �?Oo?�?fO�??O�O �O�O�O�O�O_GO,_ kO�O__�Oo_�_�_�_ �_�__oC_�_7o%o [oIoko�oo�o�_�o o�o�o3!WE g��o��o}�� ��/��S��z��� C�e�?����я��� +�m�R������s��� ����ߟ͟�E�*�i� �]�K���o������� ۯ��A�˯5�#�Y� G�}�k����	�ڿ� �����1��U�C�y� ����߿i���e���	� ��-��Qߓ�x߷�A� �ߙ��߽������)� k�P����q��� ������C�(�g��� [�I��m�������	� �� ������!WE {i������ �	SAw� ��g����/ //O/�v/�?/�/ �/�/�/�/�/?W/}/ N?�/'?�?o?�?�?�? �?�?/?OS?�?GO�? WO}OkO�O�O�OO�O +O�O__C_1_S_y_ g_�_�O�__�_�_�_ o	o?o-oOouo�_�o �_eo�o�o�o�o ;}obt+M'� �����U:�y �m�[�}����Ǐ�� �-��Q�ۏE�3�i� W�y�{���ß��)� ����A�/�e�S�u� ˟�¯������� �=�+�a�����ǯQ� ��M�˿�߿��9� {�`ϟ�)ϓρϷϥ� �������S�8�w�� k�Yߏ�}߳ߡ����� +��O���C�1�g�U� ��y����������� ��	�?�-�c�Q�������������$SER�V_MAIL  ��������OU�TPUT�����@��RV �2w�  �� �(��I��SAV�E��TOP10� 2#	 d ������ '9K]o�� ������/#/ 5/G/Y/k/}/�/�/�/ �/�/�/�/??1?C?�U?g?y?�?�?w�{Y�Pf��FZN_C�FG w����W�1GR�P 2�7t ?,B   A'@��D;� B(@��  B4�R�B21VHELL��2	w�r6 7��7�O�K%RSR �O�O�O�O�O_�O3_ _W_B_T_�_x_�_�_��_�_�_on�  ��RoKo]o+bio ��eo�b�`S�bg3b2��dul�tm�bRFHK 1
`K �o 0YTfx��� �����1�,�>��P�LLOMM �`O��QBFTOV_�ENB��+r�bO�W_REG_UI�����IMIOFW�DL����*E��WAIT���i�2�����*�TIMn���T�VA��|+���_UNIT��싖r	LCڀTRY��r��MON�_ALIAS ?5e��2 he��� !�3�E�S���v����� ��W�Я�����ï <�N�`�r���/����� ̿޿𿛿�&�8�J� ��[πϒϤ϶�a��� �����"���F�X�j� |ߎ�9߲��������� ���0�B�T���x�� �����k������� ,���P�b�t�����C� ����������(: L^	����� u� $6�Z l~��M��� �� /2/D/V/h// �/�/�/�/�//�/
? ?.?@?�/d?v?�?�? E?�?�?�?�?O�?*O <ONO`OrOO�O�O�O �O�O�O__&_8_J_ �On_�_�_�_O_�_�_ �_�_o�_4oFoXojo |o'o�o�o�o�o�o�o 0B�oSx� ��Y����� �>�P�b�t���1��� ��Ώ��򏝏�(�:� L���p���������c��ܟ� ��$�Γ�$�SMON_DEF�PROG &����N�� &*SYST�EM*+�o�����?=�RECA�LL ?}N� �( �}tpc�onn 0 >169.254.���120:1794�0 Ơ��3980� ݡ�����} �xyzrate o124=��34��̯ޯo�����&�tpdisc 05� G�H�Z�����"������Ϳ߿pςϔ� }y!*���4636K� ]��� ��%����� ����l�~ߐ�#�5�G��Y������!�:co�py frs:o�rderfil.�dat virt�:\tmpback\2���d�v����1*�mdb:*.*?�Q�6 \�����l�$�5x*�:\��4�������q�����}6*�a2�D���a��� ��)�;�����p� ���B��]�  %����[�l~����4F����/!�
��1 ���j/|/��/!md:pic�ksim_par�t1.tp�emp���/??���/ �/�/o?�?�?&,N?@G?Y?�?�?O!�2�%omay�/�?���?nO�O�O%N27OIO[O�O�O_�Ld3O�O�O h_z_�__1R�OH_Z_ �_�_o"?4?��_�_ po�o�o�?9oKo]o�o  %o�o�o�ol~ ��o5GY��� !3��h�z���� �C�U����
��/� ��ӏd�v�������?� Q�c�����+���ϟ �r������;�M�_� ���'���˯ݯn� ����%7��?��� ϣ�п�j�|ώ� !�F/W����ߟ ���U/f�xߊߝ��� 8�O�������-����Q���t����$S�NPX_ASG �2�������  0�!%�����  ?����PARAM ����� ��	��P�$� ���1�����O�FT_KB_CF�G  �#���O�PIN_SIM + ��,�����������RVNOR�DY_DO  �6�b���QSTP/_DSBv�,����SR ��� � &0�Q�'��$G�TOP_ON�_ERR����|P_TN ��� ��A�RIN�G_PRM���V�CNT_GP 2tx�.���x 	
�	� �0T��V}D� RP 1�/�E��7��� ����//1/C/ U/g/y/�/�/�/�/�/ �/�/	??-???Q?c? �?�?�?�?�?�?�?�? OO)OPOMO_OqO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_�_o!o3o EoWoio{o�o�o�o�o �o�o�o/Ah ew������ ��.�+�=�O�a�s� ��������͏��� �'�9�K�]�o����� ����ɟ۟����#� 5�G�Y���}������� ůׯ�����F�C� U�g�y���������ӿ ��	��-�?�Q�c��mPRG_COU�NTW����ENB���M��Y���_UPD 14T  
xϣ�� �/�X�S�e�wߠߛ� �߿��������0�+� =�O�x�s������ �������'�P�K� ]�o������������� ����(#5Gpk }����� � HCUg�� ������ // -/?/h/c/u/�/�/�/ �/�/�/�/??@?;? M?_?�?�?�?�?�?�? �?�?OO%O7O`O[O�mOO�O�O�O��_I�NFO 1�����P	 ��O__@_+Y@l��@I�l?Z��F_-S�̵���5Au�9�	�]�Ǝ�@���K]A�,��@� A�@�n_�D D5O�z���C�����T7��ߍ��I��Q�� 8�^NCa��ݹ. j���ּ�A���Y?SDEBUG�������@d��
`SP_�PASS��B?~kLOG �F]�  �@�X��O  ����AUD1:\Hd�NIb_MPCNm���o�o����a�o ���fSAV Qi��2Q�qa�b�E�hSV��kTEM_TIM�E 1Qg�� 0�����h��o ZwMEMBOK  ����q`�qo�� �X|&��� �_�u�"�G��W��z�����a 2[@}q��я��� /s��1�C�U�g�y� �{�����ß՟� ����/�i�e>�c� u���������ϯ�� ��)�;�M�_�q���0������\uSK�p�x���������4��@j��2,�W�A�W΀����i��Ϧ�(F��!������� ��8��%�` �-���09zm�ߑ߅��߄s���������(��@$,�P�D�t���� ����������(�:� L�^�p��������������T1SVGUNwSPD2e 'e����2MODE_LIM �vvq b2��2��Qm���ASK_OPTI�ON`�y aS_�DI+`ENB  �b�esBC2_?GRP 2ܵc|r�[R��C������BCCFG ��7| (�a� `M_VAf�w ������// /R/=/v/a/�/�/�/ �/�/�/�/??<?'? `?K?�?�?�v�;�?�? �?�?p?�?+OOOO:O sO~�O�th@�O�O�O �O�O	_�O-__=_?_ Q_�_u_�_�_�_�_�_ �_o)ooMo;oqo_o �o�o�o�o�o�o�h�0 3EW�o{i �������� �A�/�e�S�u�w��� �����я���+�� ;�a�O���s�����͟ ��ݟߟ�'��K� c�u�������5�ۯɯ ����5�G�Y�'�}� k�����ſ��տ׿� ��C�1�g�Uϋ�y� ���ϯ�����	���-� �=�?�Q߇�u߫�a� ���������;�)� K�q�_������� �����%��5�7�I� �m������������� ��!E3iW� {������� #5Sew��� ����//�=/ +/a/O/�/s/�/�/�/ �/�/?�/'??K?9? [?�?o?�?�?�?�?�? �?�?�?OGO5OkO! �O�O�O�O�OUO�O�O _1__U_g_y_G_�_ �_�_�_�_�_�_�_	o ?o-ocoQo�ouo�o�o �o�o�o�o)M ;]_q����O ���%�7��[�I� k������Ǐُ���� �!��E�3�U�W�i� ����ß���՟��� �A�/�e�S���w��� ������ѯ���+�� C�U�s�����������˿�߿���3��$�TBCSG_GR�P 2����  �3� 
 ?�  ^� p�Zϔ�~ϸϢϴ��Ϡ���$�7�>�E�_d0 �S�?3�	 HCA�"��>l�"�CS�BpVߙ�c�u߇���{B�$�>������"�Bl����)�AЎ�����G�"�;�B	�)�+�Q�G��_���A3�"�Q���T��Ѩ��@�����'� :���e���M�_��������?�ff�� ���	V3.00>V�	mt2 * 2�$��<3�G�� [ -\�  q��7�J�2>�E���C�FG !���O� R��
�r��0�0 Vd�d�u�� ����///P/ ;/t/_/�/�/�/�/�/ �/�/??:?%?^?I? �?m??�?�?�?�? O OV�p�O/OAO�?tO _O�O�O�O�O�O�O�O _(_:_L__p_[_�_ _�_�_3���_���_ ooIo7omo[o�oo �o�o�o�o�o�o3 !WEgi{�� ������-�S� A�w�e�����m�ŏ׏ ������=�+�a�O� ��s�����͟ߟ��� ��9�'�]�o����� M�����ۯɯ���� 5�#�Y�G�}�k����� ��׿ſ�����C� 1�S�U�gϝϋ��ϯ� ����	����?��W� i�{�%߫ߙ߻߽��� ���)��M�_�q�� A���������� %���5�[�I��m��� ������������! E3iW�{�� ����/? AS�w���� ���/��O/=/s/ a/�/�/�/�/�/�/? ?�/%?K?9?o?]?�? �?�?�?�?�?�?O�? !OGO5OkOYO�O}O�O �O�O�O�O_�O1__ U_C_y_g_�_�_�_�_ �_�_�_o	o+o-o?o uo��o�o�o[o�o�o �o;)_M� ���w���� �7�I�[��'���� ����ُǏ����3� !�W�E�{�i������� ��ß�����A�/� e�S�u���������� ѯ���o1�C��o�� ��s�����Ϳ��ݿ� �'�9�K�	�ρ�o� �ϓ��������Ϲ�#� �3�5�G�}�kߡߏ� �߳���������C� 1�g�U��y���� ����	���-��Q�?� a���u���%�W����� ����M;q_ ������� #%7m�� ]����/�/ !/3/i/W/�/{/�/�/ �/�/�/?�//??S? A?w?e?�?�?�?�?�? �?�?OO=OOO��gO yO�O5O�O�O�O�O�O �O_9_'_]_o_�_�_�Q_�_�_�_�_�_�^ s %`)c )f�=o)b�$TBJO�P_GRP 2"��U� / ?�)f	Ub\c�$cl��P���pJ�`��xe  � � ׸ ��`�)d �@%`tb	 �C�A��f��SC���_)eta�b33�3�f�oz=�_��CS�?���,1ru`B�;pp�gLWw�o�o?�a�u��z�<؄-r��Ͱ�u=�)eB��wC�  D�a�o�#�-�;��Bl�`2u�ff�n�)e�AЇ��w��>���ͭ�����;�{����@fff���b�]���A���������9�ˌ�X��@�o�폎���ঘ%��ɟۛ;��M���@�o���{� ���9�1�g�Y�C�Q� �����E�ϯ�ӯ� �@��կ_�y�c�q�(��пct�)f��	V3.00zcOmt2��*��yd$a)�4� F�� G9| G��v�G�/�G��� H�@H�,�H.��H�C� HYA@H�n��H�� H��� H�Y@H��`H���H��c�H��H�̿�H�nD�G� G.A G�Km Gh� G���G�x�G���G���G��:�G�ЀG��f�G���G���\��H
_��H��H���H @�H'��d�ր=L��=�#�
������)b�3o�+�)f/�?��߀f�d�RcESTPARS�hn`Rc�HR��ABLE �1%ci�)dD_�D� �@$�_�_ء_�(g0a_�	_�
�_�_ؾ�)a_��_�_�����RDI��ma�����������O�������H�����S��kc I� ����������* <N`r���� ���Hm����lb ��C,�>�P�b�� ��2�D�V�h��)NUoM  �Uma�`1` �����_CFG &+���a@U`IMEBF_TT�Ѻkc�ЎT&VER�Uj&�T#R 1'�� �8&�)b$`�! �PN  �/�/�/�/ �/	??-???Q?c?u? �?�?�?�?�?�?�?<O O)OrOMO_OuO�O�O �O�O�O�O�O__%_ 7_I_[_m__�_�_�_ �_�_�_4oo!ojoEo Womo{o�o�o�o�o�R�!_!�&@�%��MI_CHAN`'� �% .sDBGL�VL`'�%��1pE�THERAD ?U���p�/��o��o��y�1pROUmT~ !�!�t���|SNMASK�yx�#�q255.�?��=�O�a�Á�O�OLOFS_DI���ecyORQC?TRL (�+��0�ߍTΏ��'�9� K�]�o���������ɟ ۟����#�3�͏V��E�z�~�PE_DE�TAIWx��PGL�_CONFIG �.)"!��/�cell/$CID$/grp1~�@����*�<���� g�y���������P�� ��	��-�?�οc�u� �ϙϫϽ�L�^���� �)�;�M���q߃ߕ� �߹���Z�����%� 7�I�������������M}n��!�3��E�W�i��k���p�� m��������� g� DVhz��-� ���
.�R dv���;�� �//*/�N/`/r/ �/�/�/�/I/�/�/? ?&?8?�/\?n?�?�? �?�?E?�?�?�?O"O 4OFO�?jO|O�O�O�O �OSO�O�O__0_B_ �Of_x_�_�_�_�_�_�͠�User� View �}�}1234567890oo'o9oKo`]oed�`£�o���Y2�Yb_�o�o�o�o!�o�o�R3�oo������(��n4 ^#�5�G�Y�k�}�����n5�׏���� �1���R��n6Ə�� ������ӟ�D���n7z�?�Q�c�u����������n8.�����)�;�M���n�t� �lCamera�Z꯳�ſ׿������E��7�I�[� ouχϙϫϽ���ŉ  ���i���1�C� U�g�y� ϝ߯���߀����	��-�?�f�� ��]y�ߋ������� ���	��-�x�Q�c� u�������R�d��B� ��	-?Q��u �������� ��d��˰ew� ���f��/R +/=/O/a/s/�/,�� y�/�/�/�/??)? �M?_?q?�/�?�?�? �?�?�?�/d�-��?;O MO_OqO�O�O<?�O�O �O(O__%_7_I_[_ Od���O�_�_�_�_ �_o�O%o7oIo�_mo�o�o�o�o�on_�W9 So,>Pb	o s��Qo����P�(�:�ɪ	��0� u���������Ϗv� ���;�M�_�q��� ��<�N�����9�� � �$�6�H��l�~��� ۟��Ưد������ ��ۥ�Z�l�~����� ��[�ؿ���G� �2� D�V�h�z�!�[�n�� ��������� �ǿD� V�h߳όߞ߰����� �ߍϟ���}�2�D�V� h�z��3߰������ ��
��.�@�R��ߟ� F������������� ��.@��dv� ���e��Ų+U
 .@Rd�� �����//*/�  �	Y/k/ }/�/�/�/�/�/�/�/<?;   //7/ U?g?y?�?�?�?�?�? �?�?	OO-O?OQOcO uO�O�O�O�O�O�O�O __)_;_M___q_�_ �_�_�_�_�_�_oo %o7oIo[omoo�o#<�  
� (  }�M ( 	 �o �o�o�o�oC1 SUg�����:�j?: �y*� <�N��r��������� ̏������a�>� P�b�t�����ߏ��Ο ��'���(�:�L�^� ���������ʯܯ�  ��$�k�}�Z�l�~� ů����ƿؿ���C�  �2�Dϋ�h�zόϞ� ����	�����
�Q�.� @�R�d�v߈����Ͼ� ����)���*�<�N� `�߄��������� ����&�m�J�\�n� �������������3� E�"4F��j|� �����S 0BTfx��� ���//,/>/ P/���/�/�/��/ �/�/??(?o/L?^? p?�/�?�?�?�?�?�? 5?O$O6O}?ZOlO~O��O�O�O�?�p@  �B�O�O_�C�G�`���#frh:\�tpgl\rob�ots\m10i�aAS_8l.xml�Oe_w_�_�_�_�_`�_�_�_on��o >oPoboto�o�o�o�o �o�o�oo:L ^p������ � ��6�H�Z�l� ~�������Ə؏��� ��2�D�V�h�z��� ����ԟ����	� .�@�R�d�v������� ��Я�����*�<� N�`�r���������̿ ޿���&�8�J�\� nπϒϤ϶�������t�� XVA �O�+P<< )P ?���A���9�[߉� oߑ߿ߥ��������� �=�#�E�s�Y������������6�$�TPGL_OUT?PUT 1	A	A_ !�-� B�T�f�x��������� ������,>P bt�������-�!Є��2345?678901 );M_g�2� �������/ 0/B/T/f/�}p/�/ �/�/�/�/x/�/?(? :?L?^?p??~?�?�? �?�?�?�?�?$O6OHO ZOlOOO�O�O�O�O �O�O�O
_2_D_V_h_ z__�_�_�_�_�_�_ �_�_.o@oRodovo�o  o�o�o�o�o�o�o <N`r�. �������"� J�\�n�����*���ȏ@ڏ�������}рF�X�j�|�������@�#�՟�)� ( 	 ��
�@�.� d�R���v�������� Я���*��N�<�^� ��r�����̿���޿� ���J�8�n��� �8�vϨϺ͒����� ���$��
��U�g�� sߝ�w߉�����C��� ���Q�c�=��� �߁���i������ ;�M���5�����/��� ������_�q�7I ��QYk��% ����3i {���K��� �///�/e/w// �/�/�/�/�/A/�/? +?�/O?a?;?M?�?�/ ?�?�?y?�?O�?O KO]O�?aO�O-OO�O �O�O�O_oO�OG_�O 3_}_�_i_�_�_#_�_ �_o�_1oCooOoyo �_�_�o�o[o�o�o�o �o-?�ocua��������)�WGL1.XML���(��$TPOF?F_LIM ��������6�Nw_SV>�  ���P�P_MON �2��R������22�STRTC�HK 3��P��C�9�VTCOMP�ATe��T�VWV_AR 4���.i� Ə *�I����:�_DEFPROG %���%MAIN 7 TLd�T1A�3��_DISPLAY�E���Z�INST_�MSK  �� ���INUSER�叜�LCK�Q?UICKME{���Z�SCRE1������tpsc@���L�Q�P�b�_f��ST�P�RACE_CFG 5����I�	3�
?����HNL 26i�b�ѡ� ?��� )�;�M�_�q�������ITEM 27�� �%$1234567890ؿ�  =<���"�  !(�0�<��u�3�ֿ������ ��0���T�f�/ߊ�J� ��Z߀������4� >߸�b��4�F��j� ������l�������� ^������*�x��� �������6�H�l� ,��Pb��x��< � �D�(� 4���N��� �@ /dv�/$/ �~/�/��//*/�/ N/?r/2?D?�/Z?�/ �/�??�?&?�?�?~? n?�?�?�?�?0O�?�O �O�O"O�OFOXOjO�O �O:_`_r_�O~_�O_ _�_�_T_o&o�_2o �_�_�o�_�oo�o�o >o�obo�o=�oX�o h���(:L �p�B�T��x�� � �����6����l� �����k�Ə��ꏪ���� �ҟD�V����S�8��$��  ��$� ɡ{�r�
 ������үS��UD1:\߬���6�R_GRP �19Ż� 	 @{�*�<�&�\� J���n��������˿�ٺ��߯��'��?�  B�T�>�t�b� �φϼϪ�������� �:�(�^�L߂�pߒ߆��	�����4�S�CB 2:@� -�*�<�N�`�r������*�UTOR?IAL ;@�Ư��/�V_CONFIG <@�ġx��¯d��OUTPU�T =@�U���p�����������  2DVhz� R�������  2DVhz�� �����
//./ @/R/d/v/�/��/�/ �/�/�/??*?<?N? `?r?�?�?�/�?�?�? �?OO&O8OJO\OnO �O�O�?�O�O�O�O�O _"_4_F_X_j_|_�_ �O�_�_�_�_�_oo 0oBoTofoxo�o�o�_ �o�o�o�o,> Pbt���o�� ����(�:�L�^� p��������ʏ܏�  ��$�6�H�Z�l�~� ����>�P������� �(�:�L�^�p����� ������ܯ� ��$� 6�H�Z�l�~������� ůؿ���� �2�D� V�h�zόϞϰ���ӿ ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<�N�`�r�� ������������ &�8�J�\�n������� ����������"4 FXj|���� ����0BT fx������ �//,/>/P/b/t/ �/�/�/�/�/��/? ?(?:?L?^?p?�?�?�?�?�?������?�?�1�?&OɟJO \OnO�O�O�O�O�O�O �O�O_"_�/F_X_j_ |_�_�_�_�_�_�_�_ oo0oA_Tofoxo�o �o�o�o�o�o�o ,=oPbt��� ������(�9 L�^�p���������ʏ ܏� ��$�6�G�Z� l�~�������Ɵ؟� ��� �2�C�V�h�z� ������¯ԯ���
� �.�?�R�d�v����� ����п�����*� <�M�`�rτϖϨϺ� ��������&�8�I� \�n߀ߒߤ߶�����������"�4�C��$�TX_SCREE�N 1>�5;�0�}�C�� ��������u�2F t�!�3�E�W�i�{��� ������������� /��Sew��� $�H�+= O������� �V/z'/9/K/]/ o/�/��//�/�/�/ �/?#?�/�/Y?k?}? �?�?�?*?�?N?�?O�O1OCOUO�?yO�$�UALRM_MS�G ?c��p� qOFګO�O�O�O_ _6_)_;_Y___�_�_�_�_�_�ESEV � �M
f�BE�CFG @c��m�  F�@��  A:a   B�F�
 �_M�c� moo�o�o�o�o�o�o��o!/waGRPw 2A k 0F��	 Woy�@I_�BBL_NOTE� B jT���lM�h�O��,`�rDEFPRO��@%�K (%OMAINz�}%�_ ��?�*�c�N���r���������̏��{F�KEYDATA �1Cc�cpp /gF�fi�{�R��������,(���F�(�[ INST �]��  IREcCT�C�ҐND-��l�'�CHOICE��q�[EDCMD��ǯҟ�ү��� 3�E�,�i�P��������ÿ������ψ����/frh/g�ui/white�home.png�)�g�yϋϝϯπ@�instR����ϰ��*߹�  A�direc��g�yߋ� �߯�>���Q��������0��E�choicQ���u��������@�edcmd ������
��.�@���}@�arwrg�� w���������F�����  $6H��l~ ����U��  2D�hz�� ���c�
//./ @/R/�v/�/�/�/�/ �/_/�/??*?<?N? `?7�e?�?�?�?�?�? �?�/
OO.O@OROdO �?�O�O�O�O�O�OqO �O_*_<_N_`_r__ �_�_�_�_�_�__o &o8oJo\ono�_�o�o �o�o�o�o�o�o"4 FXj|��� �����0�B�T� f�x��������ҏ� �����,�>�P�b�t� �������Ο���� ���:�L�^�p�����Z/����:����ۯ�8�ɯ�(�7�,��S��POIN�T  ]\��� O�OK T ���� � NDIRECT����� CHOIC�Ew��TOUCHUP��8�\�C� ��gϤ϶ϝ������� ���4��X�j�Qߎ��m;��whitehom^���������x����poinf��R�d�v���%�Y�lookB�E���������#���indirecA�]�o�������>��choic�������'*���t?ouchup��e�w���,���arwrgL��� /&�Sew�� �<���//+/ =/�a/s/�/�/�/�/ J/�/�/??'?9?�/ ]?o?�?�?�?�?�?X? �?�?O#O5OGO�?kO }O�O�O�O�O��bO�O __1_C_U_\Oy_�_ �_�_�_�_b_�_	oo -o?oQoco�_�o�o�o �o�o�opo); M_�o����� ��~�%�7�I�[� m��������Ǐُ� z��!�3�E�W�i�{� 
�����ß՟����� �/�A�S�e�w���� ����ѯ������+� =�O�a�s���������Ϳ߿�Ϟ��}������:�@L�^�6πϒ�l�,~� ��v��������A� (�e�w�^ߛ߂߿��� �������+��O�6� s�Z��������� ��O'�9�K�]�o��� �������������� ��5GYk}� ������1 CUgy��,� ���	//�?/Q/ c/u/�/�/(/�/�/�/ �/??)?�/M?_?q? �?�?�?6?�?�?�?O O%O�?IO[OmOO�O �O�ODO�O�O�O_!_ 3_�OW_i_{_�_�_�_ @_�_�_�_oo/oAo �eowo�o�o�o�o�_ �o�o+=O�o s�����\� ��'�9�K��o��� ������ɏۏj���� #�5�G�Y��}����� ��şןf�����1� C�U�g����������� ӯ�t�	��-�?�Q� c�򯇿������Ͽ� 󿂿�)�;�M�_�q�  ϕϧϹ�������~� �%�7�I�[�m��V`����V`����߼��ݦ������,��3���W�>�{� ��t���������� ��/�A�(�e�L����� ����������  =$asRo��� ��� �'9K ]o����� ���#/5/G/Y/k/ }//�/�/�/�/�/�/ ?�/1?C?U?g?y?�? ?�?�?�?�?�?	O�? -O?OQOcOuO�O�O(O �O�O�O�O__�O;_ M___q_�_�_$_�_�_ �_�_oo%o�_Io[o moo�o�o2o�o�o�o �o!�oEWi{ �������� �/�6S�e�w����� ����N������+� =�̏a�s��������� J�ߟ���'�9�K� ڟo���������ɯX� ����#�5�G�֯k� }�������ſ׿f��� ��1�C�U��yϋ� �ϯ�����b���	�� -�?�Q�c��χߙ߫� ������p���)�;� M�_��߃������h�����p����p����,�>��`�r�L�,^��V ����������!E W>{b���� ���/S: w�p����� //+/=/O/a/p�/ �/�/�/�/�/�/�/? '?9?K?]?o?�/�?�? �?�?�?�?|?O#O5O GOYOkO}OO�O�O�O �O�O�O�O_1_C_U_ g_y__�_�_�_�_�_ �_	o�_-o?oQocouo �oo�o�o�o�o�o �o);M_q�� $������� 7�I�[�m���� ��� Ǐُ����!��E� W�i�{�������ß՟ �����/���S�e� w�������<�ѯ��� ��+���O�a�s��� ������J�߿��� '�9�ȿ]�oρϓϥ� ��F��������#�5� G���k�}ߏߡ߳��� T�������1�C��� g�y��������b� ��	��-�?�Q���u� ����������^���@);M_6�a��6������������, ��7[mT �x�����/ !//E/,/i/{/b/�/ �/�/�/�/�/�/?? A?S?2�w?�?�?�?�? �?���?OO+O=OOO aO�?�O�O�O�O�O�O nO__'_9_K_]_�O �_�_�_�_�_�_�_|_ o#o5oGoYoko�_�o �o�o�o�o�oxo 1CUgy�� ������-�?� Q�c�u��������Ϗ �����)�;�M�_� q��������˟ݟ� ���%�7�I�[�m�� ��h?��ǯٯ���� �3�E�W�i�{����� .�ÿտ����Ϭ� A�S�e�wωϛ�*Ͽ� ��������+ߺ�O� a�s߅ߗߩ�8����� ����'��K�]�o� �����F������� �#�5���Y�k�}��� ����B������� 1C��gy��� �P��	-? �cu�����ڦ���������/-�@/R/,&,>?�/6?�/�/ �/�/�/?�/%?7?? [?B??�?x?�?�?�? �?�?O�?3OOWOiO PO�OtO�O�O���O�O __/_A_Pe_w_�_ �_�_�_�_`_�_oo +o=oOo�_so�o�o�o �o�o\o�o'9 K]�o����� �j��#�5�G�Y� �}�������ŏ׏� x���1�C�U�g��� ��������ӟ�t�	� �-�?�Q�c�u���� ����ϯ�󯂯�)� ;�M�_�q� ������� ˿ݿ���O%�7�I� [�m�φ��ϵ����� ����ߞ�3�E�W�i� {ߍ�߱��������� ��/�A�S�e�w�� ��*���������� ��=�O�a�s�����&� ��������'�� K]o���4� ���#�GY k}���B�� �//1/�U/g/y/ �/�/�/>/�/�/�/	?�?-???�A;�>����j?|? �=f?�?�?�6,�O�? �OO�?;OMO4OqOXO �O�O�O�O�O�O_�O %__I_[_B__f_�_ �_�_�_�_�_�_!o3o �Woio{o�o�o�o�/ �o�o�o/A�o ew����N� ���+�=��a�s� ��������͏\��� �'�9�K�ڏo����� ����ɟX�����#� 5�G�Y��}������� ůׯf�����1�C� U��y���������ӿ �t�	��-�?�Q�c� �ϙϫϽ�����p� ��)�;�M�_�q�Ho �ߧ߹���������� %�7�I�[�m���� �����������!�3� E�W�i�{�
������� ��������/AS ew����� ��+=Oas ��&����/ /�9/K/]/o/�/�/ "/�/�/�/�/�/?#? �/G?Y?k?}?�?�?0? �?�?�?�?OO�?CO�UOgOyO�O�O�O����K�������O�O�M�O _2_V,oc_o�_n_�_�_ �_�_�_oo�_;o"o _oqoXo�o|o�o�o�o �o�o�o7I0m T�������� �!�0OE�W�i�{��� ����@�Տ����� /���S�e�w������� <�џ�����+�=� ̟a�s���������J� ߯���'�9�ȯ]� o���������ɿX�� ���#�5�G�ֿk�}� �ϡϳ���T������ �1�C�U���yߋߝ� ������b���	��-� ?�Q���u����� ������)�;�M� _�f������������ ��~�%7I[m ��������z !3EWi{
 �������/ //A/S/e/w//�/�/ �/�/�/�/?�/+?=? O?a?s?�??�?�?�? �?�?O�?'O9OKO]O oO�O�O"O�O�O�O�O �O_�O5_G_Y_k_}_ �__�_�_�_�_�_o�o�$UI_IN�USER  ����@a��   o$o_�MENHIST �1D@e � ( M`���)/SOFTP�ART/GENL�INK?curr�ent=edit�page,MAIN,1_o�o�o�o�_*�o�n"q1�oVh z�-?r2E������o�wmenu�b142�\�n�Ȁ����P(%�7�53L�M_@���	��]�-���n-BCKEDT-ُi�{����<.��mOMAYK��8���� �'�����7؏j�|������Q���P�a��ïկ�����/� ��T�f�x� ������=�ҿ���� �,ϻ�P�b�tφϘ� �ϼ�K�������(� :���^�p߂ߔߦ߸� G����� ��$�6�H� ��l�~�����ﱯ ����� �2�D�V�Y� z�����������c��� 
.@R��v� �����q *<N`���� ���m//&/8/ J/\/n/��/�/�/�/ �/�/���/"?4?F?X? j?|?/�?�?�?�?�? �?�?O0OBOTOfOxO O�O�O�O�O�O�O_ �O,_>_P_b_t_�__ �_�_�_�_�_o�_o :oLo^opo�o�o#o�o �o�o�o �/�oH Zl~���o�� ��� ��D�V�h� z�������?�ԏ��� 
��.���R�d�v��� ����;�П����� *�<�˟`�r������� ��I�ޯ���&�8��#{�$UI_PA�NEDATA 1�F���i��  	�}�  FRH/VI�SION/VRF�RMN.STM?�_imageon�ly=1&_fi�ltershow�n=0��ed=1� &_colum�ns=4��ont�=24&_p��=�wholedev�E�!v)  rim��  z�(�:�L� ^�pς�鿔ϸϟ��� �� ����6��Z�l� Sߐ�wߴ��߭���!v�� � 
��  ��"�f�rh/cgtp/�flexܰ.st�m?_width���height=�10��ܰice=�TP2&_linOes=3����1ϵ/doubܰ2���ual���$����� ����/���S�:�w� ��p����������� ��+OaH���� 
�3p��� i������% xI��m��� �.���!//E/ W/>/{/b/�/�/�/�/@�/�/�/?/?�I6 k�fk?}?�?�?�?�? ?�?\OO1OCOUO gO�?�O�O�O�O�O�O �O�O__?_&_c_u_ \_�_�_�_�_B?T?o o)o;oMo_o�_�o�? �o�o�o�o�ozo 7[B�x� ������3�E� ,�i��_�_����ÏՏ ���L��/��oS�e� w��������џ���� ��+��O�a�H��� l�������߯Ư�v� ��F�K�]�o������� ��ɿ<�����#�5� GϮ�k�}�dϡψ��� �Ͼ�������C�U� <�y�`ߝ߯�"�4��� ��	��-�?��c�ֿ �����������Z� ���;�"�_�q�X��� |�����������%I�����T������){� �8J\n��� �����/�4/ /X/j/Q/�/u/�/�/�/�/x������$U�I_POSTYP�E  ��?� 	 �/K?�2QUICKME/N  );8?N?�0RESTORE� 1G���  �*defaultx��  OUBLE~�=PRIM�?�mmenupa�ge,1422,�1�?)O;OMO_ODe�ditBMAIN O�O�O�O�O E�O�O __/_A_�1�/R_d_ �O�_�_�_�_�_�_�_ o/oAoSoeoo�o�o �o�o�o|_�o�oto =Oas�(�� �����'�9�K� ]�o�|������ۏ ����#�ƏG�Y�k� }���2���şן��� �����,���P�y��� ������d����	�� -�ЯQ�c�u�����S=oSCREi0?n=u1sc�0Wu2ڴ3ڴ4ڴU5ڴ6ڴ7ڴ8ڱTAT%=� x}3��:USER��L��Ӵksܳm�3m�U4m�5m�6m�7m��8m�0NDO_CFG H);d c�0PD�W��?None\2N��_INFO 1Ij���{00%�� �x�
�K�.�o߁�d� �߷ߚ��߾�������5�G�*�k�R<��OFFSET L)9�x�@��0H����� ������(�U�L�^� ��b������������� $6��~?�p�
����UFR+AM�0@������RTOL_ABRqT���ENB~ GRP 1M�9�z1Cz  A� ec��cu��� ���h0U/��~MSK  2��N�%����%Rs/ _EVN�2$�ƈ&��2N��
 h��U�EV!td:�\event_u�ser\w/� C7��/�B�F<�!SP��!�'spotw�eld=!C6 ????�0b$!b/�/ �?�?�7!�?�?�?O AO�?�?wO"O�OFOXO jO�O�O_�O�O�OO_ >_s__0_f_�_�_�_ �_�_o�_9oKo�_o��o,o�oPobj�&WR�K 2OXɶ8�o	 �o@R- v�c����� ��*��N�`�;��� ��q���̏��ݏ����$VARS_C�ONFI��P�� �FP@���CCRG��S��Z�@�9�D�B�BH��p����C����їϑ?��U�MRvK2Y��)�B�	��C�X�1:� SC130EFG2 *3�7�@���Y�ch �5B�����A@��CȐ� �����9���@ȯ���������ӑ��	�Z��� B���u���z� ���᯾����Ϳ� �*��'�`Ϸ�Aϖπ�ϓ�������X�TCCc�ZR�4��4pa��'�GF,��!�[�� �a 23�45678901`q�y�'9�n���n߀�ߘ#����j�����B��Ӗ ��ϑ:�o=L{��!p� � p��ia/[�ߤԆ�� ��������)�;�(� :�q��p������� ����%�I�[�H ���{��������"�>S�SELEC�$!�?�AVIA_W-O�`\T)_ff,		�= �;G�P �R'	��RTSYNCSE��j��n�eWIN?URL ?u��R���� /�/"�ISIONTwMOU�/ �*%�c�]S۳�S���@/� FR�:\,#\DATA�s?MЄ� MC�k&LOGx/   oUD1k&EX�/���' B@ ����"�!DE�SKTOP-MC6FJ6K�/�#?�%?�le � n6  ����f<�"�� -�N5K��   =�̡�w1��t0� �(TRAIN�/H҆2�b�d�3pw5{4 G#`�"'(��^]� (���9M��O O+O=OOO�OsO�O�O��O�O�O�O�O_$(S?TAT _'� � z�b_t_�_�h$�_�_�'%_GES#`]���0 �
���R��WHOMINV a/S۾�`�b"����C�ז&�WJ�MPERR 2b]�
  =�jho ^l��o�o�o�o�o�o �o.<m`r��S_� REV c\O^#�LEX�Td7���1-e�_VMPHASE  j�r��&�OFFo_ENB  \��	P2R$eSۿ�N��c|3�@�:�`Q�u���?s33�4�1K�g�']g��t�g��&�S`hWm���3�\B�c��4C�*�����&��*�Y�B��p��1��/�7k� B��a������<�	���
��� ٞ�o��,������5ǟ������j�Ϸ*��\81��_�
A/���;�M��`����O�)����� S�4�0�3��o�����[�m��������z+�CT6�<�))#X����:T�!��i����M��r/�CV�X�3�&��4�*��<C�k�}�S�M������X��^����+��~���ڿ	���O�-Od+P�kC��u�g�%�;ρ�v�^A� 
*C/嬇v���ɿ���A���MCK�߬�_�Y�K�	���e�Z�^CP�%C�p��H��#��hJ�]ݤҫ�Ϝ���M�C�b��CO��G]���+0��B�T�3� )�����C�8�X���߄�� [��� �����3���i�^� p������������  /�!S�Hw����� y������+ =2a�_q���ÅTD_FIL�TES`i�[ ����P��<//'/ 9/K/]/o/�/�/�/6 ��/�/�/??,?>?�P?b?t?�YSHIF�TMENU 1jWm<�|%��?�t �?�?O�?�?EOO.O {OROdO�O�O�O�O�O��O�O/__	LIVE/SNAP#Svsfliv�~�A_��PION� &�U^PdRmenuz___�_�_�r�5jG�kΉ��9MOG�ml�~�złZDd�m��a<ۀ �P��$WAITDINEND  �U���#bxfOK-��oO�UT�o�hS�o�iT�IM�e���lG o}�o2{�oz�oz<�o�hRELE�.�f�hTM^{d�xc_ACTWP-���h�_DATA n�΅�%�_B��6�rR�DIS�P�~�$�XVRao9n��$ZABC_GR�P 1p[k ,�2J��=Qa�pVSPT q9m����
�Z�_��Z�)�?�އDCSCHb`r#�����IPbs[o!۟����؊MPCF_G +1t�����0�� �O����u����p�� 	?���o`��  ?������{��4���c���G�4�)6C����D5Oz��ٯC��?�����<� ��>�%��6��?��u=�@p�����2?�k��1�?��Σ���4/6�u�ޤy��ꠐ>
�����������𤯎�˿ �� 8�^NC�a�ݹ. j��ּ�A���8�h����.~:��1���ڹ���&� � 2�H�Vπ˶�ȯگ�A0���� �`v�����_CYLIND��w(� ��? ,(  *E�V���B��fߣߊ�  ��������?� ��D� +�=�z�ߞ����� ���g���@�'���0v����̞�2x �� �=���?��	@��-=��`��z�A��SPHER/E 2y%���� *����X�kF X��|��� �///ewT/� x/_/q/�/��/�/�/6��ZZ�v �f