��  	c4�A��*SYST�EM*��V9.1�0214 8/�21/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA�RA�  �  �AIO_C�NV� l� R�AC�LO�MO�D_TYP@FI�R�HAL�>#I�N_OU�FAC�� gINTERC�EPfBI�IZ�@!LRM_RE�CO"  � A�LM�"ENB���&ON�!� MDG�/ 0 $DEBUG1A�"d
�$3AO� ."��!�_IF� � 
$ENABL@QC#� P dC#U5K�!MA�B �"��
� OG�f 0COURR_D1P $Q3GLIN@S1I4$C$�AUSOd�APPINFOEQ/� �L A �?1�5/ H ��79EQUIP� 2�0NAM�� ��2_OVR��$VERSI� ���0COU�PLE,   �$�!PPV1CESH C G1�!�PR0��2	 � $�SOFT�T_I�DBTOTAL_�EQ� Q1]@NO�`BU SPI_IN�DE]uEXBSC_REEN_�4B7SIG�0O%K�W@PK_FI0	$THKY�GoPANEhD � �DUMMY1dH�D�!U4 Q!RG1�R�
 � $TIT1d ��� �7Td7T� 7TP7T5�5V65V75V85V95W05W>W�A7URWQT7UfW1pW1zW1�W�1�W 6P!SBN�_CF�!�0�$!J� ; 
2�1_�CMNT�$F�LAGS]�CH�E"$Nb_OP�T�2p�(CEL�LSETUP 7 `�0HO�0 �PRZ1%{cMAC{RO�bREPR�hD0D+t@��b{�e[HM MN�B
1^�UTOB U��0 9DoEVIC4STI�0��� P@13��`B�Qdf"VAL�#IS�P_UNI�#p_�DOv7IyFR_F�@K%D13�;A�c�C_WA?t�a�z�OFF_@N�DEL�xLF0q�A�q�r?q�p�C?�`�A�E�C#�s�A�TB�t�d�MO<� �sE � [�M�s��2�REV��BILF��1XI�� %�R  �� OD}`j�$NO`M�+��b�x�/�"u�� �����!X�@Dd� p E RD_�Eb��$FSS�B�&W`KBD_S�E2uAG� G�2B "_��B�� V�tp:5`ׁQC ��a�_EDu � �S C2��`S�p��4%$l �t$O�P�@QB�qy�_OqK���0, P_C� �y��dh�U �`LACI�!�a���� Fq�COMM� �0$D��ϑ�@�pX��OR� BIGALLOW� (KD2�2�@VAR5�d!�A�B e`BL[@S �C ,KJqM�H`S�p�Z@M_O]z��w�CFd X�0�GR@��M�N�FLI���;@UI�RE�84�"� SW�IT=$/0_No`S��"CFd0M�{ �#PEED��@!�%`���p3`J3t	V�&$E�..p`|L��ELBOF�  �m��m�p/0��C	P�� F�B����1x��r@1J1E_y_T>!Բ�`��gt���G� �0WARNMxp�d�%`�V`NST� C�OR-rFLT�R�TRAT T|�`� $ACCq�M�� R�r$OR�I�.&ӧRT�S�Fg�0CHGV0I��p�T��PA�I�{�T�!��� � �#@a����HDR�B��2�BJP; �C��3�4�U5�6�7�8��9>���x@�2 ]@� TRQ��$%fh��ր����_U�������Oc <�� ����Ȩ3�2��L�LECM�-�MULTIV4�"$��A
2>q�CHILD>�
1���z@T_1b ; 4� STY2�b4�=@�)24����@�� |9$��T�A�I`�E��eT�O���E��EXT����ᗑ�B��22Q�0>��@��01b.'��B ��A�K�  �"K�/%�a��@R���?s��=�O�!M���;A�֗�M�� 	��  =�I�" �L�0[�� R�pA��$JOBB������`���IGI�# d Ӏ����R�-'r��A�ҧ��_M��b$� tӀFL6�BN9G�A��TBA� ϑ �!��
/1�À�0���R0�P/p ����%�|��Bq@4W�
2JW�_RH�ECZJZ�_zJ?�D/5C�	�ӧ��@�����Rd&� !����ǯ�rGӨg@�NHANC��$LG/��a2qӐ� ـ@�B�A�p� ���aR�`�>$x��?#DB�f?#RA�c?#AZt@��(.�����`FCT�����_F࠳`�S	M��!I�+lA�%`  �` ���$/�/�� ��[�a��M�0\�ؿ`��أHK��AEPs@͐�!�"W��N� �S'�I��' � . II��2�(>p�STD_C�t�1\Q��USTڒU�)#�0U[�%?I-O1��� _Up�q��* \��=�AO�RzsBp;�]��`O,6  RSY�G�0�q >EUp��H`G�� {@]��DBPXWORK��+��$SKP9_�pAqfau�0��TR�p , ��=�`����Z m�OD3��a _C"�;b�C� �GPL:c�a�tő"S�D��G�Bb`����P�.� )�DB�!�-|B AP=R��
 �DJa3��. /�u����� �LUY/b_tS���0�_���PCr�1�_�TENEG��]� 2�_�S6PR�E.��R3H {$C��.$Lc�/$USނz )kIN�E�7A_D1%�ROyp�������qbc�7 T@zfPA���R�ETURNxb�M�MR"U��I�CR�G`EWM�0�SIGNZ�A ���e�� 0$P'�g1$P� m�2�`B��`tm�pDIp� �'�Bd.a	r�GO_AW ���0ؑ�B1m@CSd�(�C%YI�4���`1wsqTu�|t2vz2�vN��}��E]sDEVI�S` 5 P M$��RB��I�wyPk��vI_BY����p�TQ�tHND=G�Q6 H4��1��w��$DSBL C��O��vG@��SP_qL��7/�F@]�d�3FB���FERa8�����t]s���8> pi�T1?���MCS솠��FD ���[2H� W ��EE���%F��Żt�SLAd��09  ��INP^��]�`�|]q��:P +8�S��0x�^���^���FI�2��������A	AWl���N�TV�㜒V~���SKI�#TE����a����T1J_�#;2_��PD�SAF�T�_�SV�EXCLUT�῰�D6@Ll ��Yք��3�HI_yV
0\2PPLY�@�0«�G�����_ML�%��pVRFY_t�C��M��IOC�UC_� ���O��p��LS�`V�&T4��A1��s���@P�dE&�gp�AU��NFT�u��uZ��pm�ACHD�O���^����AFC CPl��T�D�4P~�� �� ;��P@T�ѡ0,@ '��I���N��=�' <Y���T��?�q ���{�SGN��=;
$�`�a>a R0I�3�g@ _BM�_B>]�ANNUN�P~� �ÅuC.@�`/���ɢ�� �����2EF�C@I�R>p�$F���4OT�`{�&T�D�(RQ<�#QmJ�Mb�NI�R?��4һr6�A��R�DAYCLOAD�tT-�'S�5#Q�EFF_WAXI��@�PQ�O3O�йS�@_RT;RQ��A D1�	`���Q,@ ��EVp�Ӓ���@�0}�0X��{��MP�E{� BV�����L$s��DU�`����B�CAB��C���PN�S"�+0ID�WR����V!� V�wV_8���V �DI� �4D� 1$V�`SEm�TQj}�`'���D�^E_nѶ$�VE� � SW���[a�����A��OH��)�P�P��%�IR�1B u@p�&���b����]� w3W�O � W��vM����C�0��cp��RQD�WF�MSw0��AXx,���$�LIFE�@����-Q��N��H����Co���CB0LqN]a���3OV0HEQ�'SUP�T����@_oS�1_��Gq
�Z�
W�
B1��#��@�k2XZ_ LQ+Y2�C9`T_@``���N�����J�! �>�_� ��F� �4�E `�pCACH8,�\�]SIZ(T ��bN�UFFI� ���@(T��2'S6#Q�1DMp0��F 8��KEYI7MAG�cTM,aV#���a�^�hB1�OC'VIE�aG�2� �L��H���?� 	R��D� PH���ST'�!C"D�K$�PK$-�K$��K EMAILK�u`[��0��/FAUL�RI�2sc�C� COU�0iA�0�T`�1J< �$�#�S�m�ITW�BUFp��p�t��0�0n B�$�tCු���"�3� SAV -5�"����H7@@���P44�
`�N�_0� 5LЉ9OTgb+����P�P�:���7AXC����X� T�a3�_G��
m@YN_\N� K <\�D�uTPb�M�M8�H 5TL�F~`$�`��DIزE�@`�aILY���G1��&G��Da:AF����baMa�`A�#�3C_^`��`Knd�@^DQ�Rp��E�(ADSP�6BPC�KIM:3�C�A��A��U�Gd meڠ� IP��C7�3��DTH���B��T�aa�CHSEC�CBSC	�"�PV���Z�P��3�Tp��NVk�G �S�T�F� F���0ad�C5@�1aSC���u�CMER��QF�BCMP��~@ETn;� N�FU� �DU� ́�`���CaD�IYP�0�#m��`SNOu�=�O���p�zbL�xds�P�zbC""��e
��2�!uc|�0� PH *�aL��_c�q�1f��,� '��dD��f"��f-��fP���f��f7�i8�i�9�j���hz1z1�z1(z15z1Bz1�Oz1\z1iz2wz2T{z2z2(z25zU2Bz2Oz2\z2iz�3wz3z3{z3�(z35z3Bz3Oz3�\z3iz4wr�EX	T��=�QB\h@%�@�e@C��e�0F{DR��RT� �VW��2�򁑇R��R�EM��Fq��OV�M�C��A��TRO�V��DT80КMX�ߜIN��: Ϛ��IND���
�F@�0@G�1d�ِ9 ��9D��ِRIV԰&���GEAR�AIO��K��$�N5@���������� %�Z_MsCM� ���Fe ;UR3bS ,�a1�? 9 P?\���?�E,� ���1`v�T���5P�1��RI^e����#ETUP2_ gU -��#TDGP0��$Ti��Z�T�qa��"BACBV T(D��"eD)_J%�ýc0@ѰIFI:�0@`��`�Ь�PT��L{UI6$W �� (� URt�1@�2�MA�P� ����I��$�(�Sܰ?x4�J�b@CO|0�3VRT|$���x$SHO�����#ASSjP�1(IPQ�BG_����s���s��(s��5sFO�RC�"7��DAT�A��X�"FUס1t:B��2:ALOG����Y |*�NA�V�0�(�X���S�"&$VI�SI[�.BSC�4SQE�t�7�VB�Or���Bò�A�Z��$PO,�IE���FMR2s�Z ��i`f⁑s@ �օ�������ǖ� ��ʠ�_wqX���IT_ֱSd��ME�j�|��DGCLF;�DG�DYd�LD�H�5�
?�ѡMcp8#[���� T�F9S�07$\ P2���|sC�0$EX_������1�0�PE��3��5��G�Q��]� ��0bSW5O>��DEBUG��]񦥕GRc��U�SB�KU`O1�p  PO�Ј�t�"`tG�t�Ms�LOO�3��SM�E<2|���& _E ^ ���TERM��_���� ORISA��`<��cp�SM_`@]�B��a������ b���~�UP"c� -�D�^(���f �_>�Gk
}�ELT�O�!>B�PFIG�f?AנS�`b`�$UFRfB$`{`�� Ne�OT�ƾPTAiP���NSTT@PAT^Qi�OPTHJ&aL`E9 8d2U`�ARTU0�p� U1�">ARELAc1SHFTPR?A�3__�R/`Ic ) $8�b.႐S��S�2SHId+�Uz�b O1AYLO.P �1 A��j����e[PERV p� $��T@A��Ȱ+%���ȰRC��eASY1M3A�e?AWJ�$�� �E$�/[)�OaU�$T@ A3��&IP�S��Q�ORT@MF��/����d���t��� �16�HOs���e �˶sЖi`OC���$OP^��A�cv�#��a�i@��R0�R�S"OU�Se�R�5m8K���e$PWR]�IM�5"R_H3(*� �?AUD$�kSV�oc1SDfH�$HzdE!@ADDRC�H��G7A,A%A"��p@F��ag H2�S �PFѝ�dE��dEsdE�(sSE��H��`HSvY`MN�hW�`@0��"QebaOL/S�W�{0R�\f��ACR�O����ND_C�/Szb��4�QROU	P�S2_��
Ғ�11�q��:S�DY3 DY ��EXpDY(pDY�����AC���SAVED�?W�SOUG�C��i3 $��@0_D)���j«BPRM_
��~�HTTP_z`H��aj (;`OBJ�B�%B��$C�LE��0a�`k � Q4��6�_�T���XbS0�3��KRL~�9HITCOU����G�LS�j0Xbb�$�0f�j0ʷk0SS���d�JQUERY_F�LA�C_ _WEBwSOCI��HWcqԛ+�l_@� IN'CPU�R*�Ovma ��K�0pzD/q�D/qǂ��IOLN��m� 82�R��i�$�SL��$INP7UT_��$�0~x�Py� mZpSL�P+�nep{�u�t�B#�uB"NAIO�PF�_AS��o��$(��B��qN�Y��2���ksM�ts�HY�B�5���A�pUOP��p `�pS�C��� %���,�}��0P�3�0�s���,������IP�_ME\��q X��pIP,@�Rւ_NP��`*�G2B��O��BSP���P���#BG�Q�-�M<!�gr l �TA�3`As�TI���%� ���_�OPS^�BU��ID�Ўbs���x0`��;a-���� s�r"?�r�S��pNҘ���ӕ�IRCA_C}N� t �Jim�pCY�@EA� �C��q��31�#��@xz"���!DAY_����NTVA����u�p�r#��u�SCA�Fu�CLO᎑j����@��u��ڔ$��N_R0Cβ򐎒c�6�v�r��^3%���'b������Pi��� 2Gu �����w��8\�'b\�LAB�z�\�Ѐ�UNIбn�	 ITYl�.�0E���R; G���x�r�R�_URLЀ$A�AEN|�k�*��0�C�T�AT_U#� �iJp��yр$_%E�pRk�.��A�S��q8�J�aC�FL���K��P
W�r�
�wUJR�%z �J`AF��(����D£�$J7S%�J8B��7&�h�����7���8�ɭ�APHI��Q����D��J�7J8"�L_K�E��  �K�QpLMܑ { �<٠XR�p$p�WATCH_VA�Ax�ű#fFIEL�b"Cy��2Ҳ�| 
�b�V�G-1��CTܰ�������LGɳ�}� !�LG_SIZRdv��հ�X���p��FD��I�� �ة�����������d3 ��V��V��pV��V���V�K!G�� _� _�CM�������F �!�����А4(�Ѡ���������p��� �I��
�����������RSU� � (.p�LNԢ��"~_��`DE��E�r!�s���S��r0L���DAU���EA�PQp44���GqH52X��pBOOYA?� C�ʀ�IT�c��� �RE4�SCR��|c��D�PKr,QMARGI�q�;�v�S4e$�d�qS8c�rWC�qܕ��JGM�MN3CH���qFN(Ҟ1K����	UF��n�FWD�HLSTP�
V����,���RS?H� ��C�~"�� w�U�Q�v���d��G�	PPO��"2�� ��	E]X�TUI�I;� ��;�8bZ#�Z#� ���R��P# #9N�A�3ANA�rA1���AI���D�� �D�CSf�lC�#zC�"O��(O�'SK�2�(S�(ZIGN�Ў��0���4��$DEA|�LL"�
��q���Ѐ4�м�T��$�׳��r
���n2�A�B��۠lp*s�A��+S1�52�53�1.�8"� �Ђ �Jk�0�$�u�t���Q�e����:FSTe�R��Y�B\A �$EkFCkK���PzFp�F��#�у Lp #�n�8����Co`��d��P�Dtm�}#_ � �Pt��P���$ S�MCt��� �J`CLDP|e� �TRQLI��"�PY>TFL%�iR�Q�rS��D��rWpLD8rU\TrUORG(�v��R��RESERV 2t�T>s�TIr /Sv�?� � 	[Uv�MTrUSVd�PP^�	��Q+d3fRCLMCAd�_�_SiTp3a|�OMDBG�qͰ�?��$DEBUGMCAS&�_�P���Uu�T� |�E�����MFRQV��� � ��HRS�_RU�q�A'�A<5��FREQ�����$� ��OVER�t���F��P�EFI��%�A(��ar���c�T� \��q��$U@%�3?`��PS�0C�	sC��BcN��sSc�Uݐ�a?( 	�{�MISCuŊ Yd}�ARQA�	�3TBN �� �m!��AX �-��.�E�XCES벽��rM��̱����r ľ���rSC@ � 	H"�	�_S��8���(,�>�.PKɴ��r���N �eB_��FLI�C�DB QUIR-E�MO��O�pv��QL�@Mȵ� @P��E����Ab�a#ND��q�ހ�{�r���؄�D���INAsUT4��RSM�����+0N$bn�j�PwSTḺ� 4٠7LOCFRI��E;EX�ANG�"�qn�aODA�e��p1|����MF��� Cv7I�BA �Eq�o�fgSUP�EwqFX;��IGG � �`�Cn�(�C��D a�br\B��^@ɨ^@ئ`���P��7�qTIv�Ȼ��Po�M+��b� Mt9�MD6���)D�� O�XaL�H���O�GDIA��P�>�WiPO��1�O�D��)/��t�)`ހ� m�C�U��V��#`�qՁOr\_�`y�� ���0CC��`rr�� ȡP �J���P��KqE�^���-$B+p��@ND2ZbZ�P��2_TX�DXTR�A�#|�lb�E�LOľ�ހ�k���� ���u�ǲ�ƪ�%�R�R2�u�� .�����A0a d$OCALI�o�G�!:��2�0RIN����w<$R��SW0_d�,�lcABCJ�D_�Jb����pC�_J3:W�
Q�1SP�Т��pPQ�x�3w�̱�@
�p��Jlc���R(a�Ou1IMl`�rCS�KP_Z�Ի��#��J���rQ��������_AZ/b��I�E�LZ1��ZaOCMP0��q�q��RT�at�Ƥ�1��В��1���{ ��Z��SMG�Y'�zdJGPSCyLN�
�SPH_0��p7��㓰�p��R'TER+���� ��)_� Q6@A\ SC��r'�DI_���23�U��DF{�H�L�WN�VELPQIN8�Bf q�_BL� �ry��ѳqJi�~������MECH�2lbwqIN
�q���ǲ��]Ҳq ��@_�p ������/��`�􆂛��?�ՀDHN�~�����0$V������{!$��'qrA��$O1.PR������H �$BEL�Z��g�_ACCE�� �la� IR�C_(��a�PNT<�q;C$PSN�CRL{���XS��� ?�� �G��	�3�ؠQ�_�1lIpO"u�p�_MGscDDl(�rFW3P�(�����}DE��PPABN�RO��EE_�1�PP���1�a���{�$OUSE_���#P+pCTR�$Y�~ .a- �AYN�pAm 6&��f�6!M�aұ�"fqOk�
c$INC��������'���ENC�L��r��,�� INCBI��%�)���NTi��NT�23_L�r�#LO]�r09pI\��6�R���p���0����C<���&MOSIq���߰O!s�rPERCGH  ��7q� y7 ��3�2zd�o�g� %&N��A��5L $�ӻ����%��:F�36TRK��AAY ���3��HA�WELC�pz暁�"�`MOM}"�����P̰����0cC���DU��D�S_BCKLSH_C��E�`X68p>#��s�C�"ZM!�CLALM�$�a�@ 5U�CHK���Z�GLRTY��A��$��Qr'�_f�M4_UM�c��VC�cz��SpLMTt�_Lj b�Tv��WE�]�P�[�P���U��нc�2 d�8P	C�1�8H��&�p�U�CMC��z~CN�_	�N��f��SF��9V "��'�Ta���eXhCAT�^SHf�	�~�&yQ�A�&`����ɗ�mPA�T&�"_P�UrC_�����OFm0��_CqtbUJG0J�d�esW�OGrg�TORQU ��K3�hI��c2��r_W�EHD��m�t^�uTd�uI�{I
�Id�F0��q��I���vVEC� 0����j�1p�pn��0�v�JRKp�X������DB��M��:��M��_DL^�2GRV�t�^�d�ՁH_��Ӄ"�CcOS/�|�/�LN�� R�s�Y�^ T���T�&���~�D�ЅZM�c6ՁMY[�Θ;�I�C���THET0#5NK�23d�X\�CB��CBXC��AS��C�&�Q�^Q��SqB^o�)�GTS���C{�Kq��:s�祪��$DU_P�7ʢP��٧��Q�1_4cVqNE��KoT��-�< �A�:�C�8!�,�,�LPH/���%�Ss���~�����@���������:�V\�QVQ�N t�V��V��UV��V��V��VȻVֹH\�u�{�s��aT�Ȑ�H��H��H��UHȻHֹOM�O\��O�r�O��O��O���O��O��OȻO��F�>���~���O��SPBALANC�E_ޑ��LE��H_�SP��o���~�|�ҍ�PFULC��`��⍕��1����UTO_ZPbUT13T2^�2NAQ� � ~���A�������AT	@OA��pI�NSEG�<1REqV��<0�!DIF2Ef	1���?�1�%@COB��%Q���G2�p�� LQ݄LCHWA�R�%"ABAq�E@��<0ސU!���SXUA�Pdt�3�?S�� �
u��q��%ROB�m0CR�2��ib � �C�_]rT �� x $W�EIGHR p$�M���tpIR!0IF�
!�LAGC""bS�C"��C"BIL)O1D�@?0ST� P��%P  | �`��
����
� �D!]q�  2�J4DEKBULXɠOMMY9���N+s��p$D�1�$� op �  _ �DO_� A��� <��rh��D!�0�BB: N�#_�!0D _O2P _�� %�PT� ��!�QT��� TI�CK-�T1� %j�@sNm0M�	m0R�@D!=�=�� _PROMPR#E/�? $IR�pB!phP��0"MAIڀh}!T"�_# ����^AV R�COD�wFUJ ID_��0'%�����G_SwUFF&� 49!��DO����< �GR#=�e$ �q$=�|%=�%�qe$��� ���H�_F�Iv9�#ORDfB ��36b��"B!� $ZDT�.%�0_��4 =*��L_NAs|52�DEF_IE8 52�Q4�I�S�0}3��5�IS��` ���3�O4�a"�4�abSDQ��B��4wD�pO�� LOCKE+q_#��0��1e"_ UMd%52 e$}3e$�5e$�2q"gC p%`3q$�4q"Q�F�1 |#H�^q|%52|%}3|#�GUa(8P�4H��1�� WFHEU<C� 1TE0Q��� LOMB_t_RzW0VIS=�WITYAoqOCA_FRIN�S�#SI�1�Q�Rp�W�{�W3�W�XW��[倩V��_i�!EAS�"�q�Tp@T��V4�Y5�Y6�ORMULA_I�+q�G%7� h� �7�COEFF_OW��dW���GqS �CaA���_GR�� � � $h<@��
XGTM/G�'t<E]DCA|ER���T%D$4� �  �G�LL�$@S/�_3SV�4�x$hV� q����d� � r�SETU�3MEA��D b� _�"��� � �p��  � �` �� �A�:2�sA0AD�b �Q�";��@�1@�G����RECt�!�2SK_���s� P��1_USERz�j���,�8����z�VEL>����,�����=�I0����MT8CFG���O  u��Oc�NORE�� ���-��� 4 p�s^�d�XYZ�#��������_ERR�� ��ep6 A�c\�}��Ҁ� BUFINDX1�t��PRt� H��CU\�d��1xӃ���!$������10� 1���G�r� � $S�I�`�P �ᝀVOx
����OBJE��ADJU����AY9p���DJ�O�U� 5���C!�"=��T��y���x��DIR}��������⎴�DYNb����T�R�5�R�QHB 4���OPWOR� ��,� SYSB9U*�2�SOP��$�q�U���P<@߂4�PA���6�_�2�+OPz U4�(��xt�e�IMAGo�1��q�SIM���IN`\���RGO�VRD��%���g�P i��������@ C׵d��L:@BY��� �PMGC_E0��N*�M±�1�2��sSL���� ���OVSL��S:RD#EX�1�0K�2c���a_��cǬ ��cì  mÂ�}Ȫ��C��70����Ƿ�_ZER� �*��s��� @h"���~�O/ RI���
��������T��'�L�����T`�W ATUS�p�C#_T����O�B+pYրB���3�.�0��� D�e�N�LҾ��`M��!��o��XES� ��һ҆��ò�����R�UP:��0�1PX��y�b��3ǂ� ��PG텳��$SUBA�~��AA��JMPWAIT��r�Y�LOW/�^�' CVF�vc�\�R���q�CC��R���i��IGNR_{PL�DBTBW P�1d�BW ����U*��IGL��I�c�TNLN����R�֡5B�PN�E�PE�ED��T�HADO!WW b���ES�M��b�+�P0SPD��� L��Ar�Q0m�/��{�UN �y���R��м�LY0��K��'�PH_PK��~��RETRIEӌ�i�y!0���FI�� �:������ 2���DBG�LV��LOGSIYZ��1KTy�U�sr2D8� �_TX�EM�`Cn���X A�RR.R+�CHEC9K��1��P��p�e�c�����LE�4pPA#@T��C�O�қP��p�bAR@%"���#�1'�O� 0��`ATT���x��%X ��1��UX����PL, � $��/QSWIT�CHT��aW�ASr���SLLBp���� $BArv�D
C2�BAM��h�����J5L����6�|_KN�OW����U=�A�D��`x�D��)PAYLOA��@%#�_��.'�.'Z+#L�AA�q�0LCL_ʐ !�pg"��Ӂt$˲�&F�)C�gpb*�e$�`Ib(R�ipb'{�~$B7`ʑJL���!_Jl!��֑ANDz�U�
4l"�!�(�"aPL�AL_ �`x�ѐ�����PC>�D*#E=��sJ3036� T�`�PDCK�22�C}O�p_ALPHC3��3BEБsaC?U<���b��� � ��.�$/D_1+*2U$D�pAR��H�5xFC�TIA41Iu51I6>�MOM��@=C]CJC]CWC�Bp��AD=C�FJC�FWCPUB�RbD�EJC�E�WB�@30ʑq� � � MO"L�� �T���� e$PI����3@��0'&Y��J)&YI2[I@[INS�DS�V�V�ޠ2������1�HIGo1�q�j� �Vj�q�����V�S�X���Y��q�SAMP �Я�:d�W;cq�3 �piaʐS�Œ xd��fj��0�i@Œ@ߠ�:@�e/0��H��cIN�l/0c�h�k��dq��jx�d{2{G�AMM�eSU�A��$GET�R��3�D��4҂
$60IBRt���IL�$HI:�!_����Œ�vEѐ�x1A�~�p�vLW�}�v �|�y��v�2�V�51C��CHKİ��q�x>I_`�ޔ.2 �8.1�e|�uCޔ�F{��33 �$e8 �1��I�RC�H_D����RNs�8���LE���R�����8Ѐ��MSWsFL���ASCR�G100{�. xd39 ]��gʐ=@�iq�j����PI3AVMET�HO�æ��妒AX�$���X4�p�ESRI��:d3fsR�� 5	�Q�0FWt;acI��c�(�L�;a=�OOPa֑S���a֑APP��F�� W�x�c��cRT��2�O0j�0�������DR 1�%��D���ѪNPѢRA� MG��OSV	Q��P; CURC��G�RO7���S_SA��ܴ5���NO�0C �����45��t�?6/H/ TX����zP��UϸCDOi�A�rdyes� �e�X��W��X3�/���k#���D�T� 7� ��YL$S�!
�g��S�"6A9�ǂK���!�����!_r�C���M_Wd�B��C�����?�M�� �ˇ ��21~�L�T��K�� PM&�R� !�}�R��WE�S$��L3X!EШ4 Cү4CҶ4C�W4���pAN��sf��/0X��	O�3.1Z�� P{�TW� ���M��z� w���������4@������ �C�1_Z� | v1��5�]I��JC��WC�5�6J���PJuu Q9 p�����Y �s�P��PMON�_QU?` � =8� QCOU��7QTH_�HO~�:�7HYSES�:�UE%�+�� OXǋ  ��P#ПuV�R_UN_TO����9O�R
P� P! ���C����INDE>�ROGRA��J���2C�NE_NO����IT�A��g�IwNFO��� bh��������OI���� (SLEQ��V"�U" ��A�OS�U��� 4� E�NABqҁ�PTI�ON
�ERVE��R~�Q�VGCF._� @.�J �.1V����pR����T_EDITN��� �R���K�Aj�S�qE�pNU�AUTQ�	CO�PY�A�P*�Q]�M�qN48M�PRU�TR ;N� OUC�Q$G�����RGADJ��� -hv0X_��I����(��пW�P��п�S��rN0_C�YCq��RGN�S[�s�=�LGO�Z��PNYQ_FR�EQ�BW�`�VP!S3IZn[�LAœG!p�XC�`�UCRE�p̸�[�IF@Q��NA�Ca%�$_GœS�TATUv�œy�MAILAb�1�!
�5�LAST�!�1"$EwLEM_� �\�>iFEASIl3� nbg�Z�2��>�96���`�pI����G"�Q=� ��n2ABU�0E����PV�!�6BAS�2�5�r�AU�P�PJ�g$�1�7RM�@Rh3Ł���3���P�r��!�4 ��$"S��~�	E2 2� �c���d+F�2*G �2"Э`���2VGW��DOU����r�"$P� �@�)GRID���U�BARS�WT9Ym "OTO����W� t�_�$!���B�DO��\� �s ����POR���C���CSRV� )lTVDIS�T_�P@4PFT�PPW�PPW4NYU5NY6NY7NY82Q��Fbr_�r�$VALU�3(�+4��|�Q\�� !h�^����C�!%���A�N'��R�!��T")1TOTAL_�$l06b�PW=#I�AKdREGGENIj^b��X�8`��=�� f �TR�3�"Ia_S+��g^`��AV���b��2E�#� �?�(2�� cV_�H�@DA ��`pS�_YY���a&S8�A�R �2� �IG_SE6�`R�%�_���dC_�F$C�Mm�f�wrDEh�?p�rI]�ZvsPsq!z�F��HANC&�O� pAj�"d#qINT1P��yF}���MASK��0OVR��� �<�0�!Ł�Gy����Q�E��d�OJ6�k�F�P�SLGHp�Q� \ 1�b%Z�$�3`� qS���$�qUY��y����c��ZQUs�T�E��@� (ĆaJV�Q�q#IL_Mp$�Vt2����CTQ ����0C��j��VB�CP�P_��J�Z�Mq�V1p�VU1~�2��2~�3��3~�4��4~�� �`�<�����IN�VIB0�J�7��>�U2:�2F�3:�3F�4:�4F���Y�r�U� �gP
�tP��'��;PL� TOR$�ŃIN��u�5�����T $MC_YFC�X��LC�(B��u)`M��I�s*��rC ��)�r��K�EEP_HNADED#�!e��0o�C�т�����A$�����O �d�>"��`���w��REM�����!�B�µٱ޸U�$e��HPWD  e��SBM�q�@COLLAB"��P��'a�"� IT' ��IN=O)�FCALh�
�n��� ,��FLn�>�1$SYN����M��Ccr��`UP�_DLY���r�DGELA���!�"Y ��AD �.�QSK;IPG�� �
P��aO��˂K���P_�� ���Ƕ�����#� �#�gP"�tP"ځP"�@�P"ڛP"ڨP"�9�O�J2R ���dX�0TJ#����)1����a�����a��RD�Caw�� �� R��R�!�=��-D�RGE� W3�{BFcLG�0��SW{	�-DSPC��!UM�_����2TH2N�uA��� 1ߏ  ����A[ � D���x]�0O2_PC���S��|�1Q L10_Co"8����q ��� JPٰ7��6K�+��� �.�NE���N�0��b\r�3���p�����DESIG\��JEVL1��1���k��10ٰ_DS`�K�j��`C11��� lV�������iI�AT����AS'J N$	C�
����HOME4 ���2�������� 2D����3����gy���� ��4�����P,>�5���a`s���� ��
�6�����//(&/8/V7���[/m/�/�/�/�/J'8�����/�/�/? ?2? R��S)������1���s`Y�V۰E�D�� T���4,f�3IIO��
II�0XrOe�_OPE.C&b�3��POWE�� �0�����P/�'c� �}�eB$DSB��GNAr�%c���C���Q�S232N�5� ��Z5���׀ICEUS/cS�PE���QPARI9Tq$aOPBQ��RoFLOWApTR�041b�UJsCU�@6���QUXT�q�Q�pEORFAC�DʰU `�J"SCH�Q� tV��_�@kpc�3$�`�`OM*p���A>�#�p%�UPD�<����aPT�0|uE�XЙX|S!%�FA�?��r��q�a � ���`;b K�AEL$� ��U��]B��a  2� ��S���0�	� ��${�����GRO��`*dT�(p6fD;SPBfJOG�`�C����AZ�N�������"VK�P_MIR�^a~d�MT3��cA�P%����`}t��S�p�`R��
��eBR�KHUQ�V��AXI�1  �bc�r-b��q9�7e�`BSOC�6f۰N2uDUMM�Y16O�$SV&��DE3A�CF�wK�e0�D�pcOR{ws0N�p|vFp�w[`�OV^eSF�zRU�N�s�rF�vQ�cU�FRA�zTOTLcCH�����OVlt[�[`WP�7�[c���r�?p��_�p� @>h�TINVEG@n1�OFS\�C�P�WD�q��q>qf2�eXp�TRr��1a�E_�FD�aMB_CW���B��B�*��ałˁ?�epV9Q��P�&��írGƇ�hAM��c��VP�F�!�_M`݀R_�CS�T$�����Q�3T$HBKX�Q�fm�IO�5|�&A��PPAp�����ଔ��,�&BS�DVC_DBъ0ސ�Q�B ސ7�Q������F���3��L�E���+P�`lqqU�3P`FCAB�Ѐ�2~㷀8û` ���O��UX�fSUBCP�[�-��/���P/Ѯ�ރ�bB��$HW_C��	P/ш���?�q0#��P��$UP�t	��A�TTRIh��h`C3YC��g�CAB��c�FLTR_2_FAI�3�IH��F��Ptk�CHK�_SCT6�cF_�F_�����FS�A��CH�A�}�ֱ�RղRSD���Aq�S�A&@�_T�}�.���PE)M�0��MsTò/���Pò��K�DIA�G�URAILAC4듑�M`LO"p��<Hv_�$PSNb�2� ��L��PRߐS�}�I���Cёf�	�E�FUN��*QRIN1�}�|0^���Q&�S_;`��X�����0f���P�f�CBL���.�A'�#�*�#؃DAp��h�.�'�L�DyP`p����Ca�����TI�°���P�$CE_RIA�a�BAF��P�AX��~���T2}�C�S��؁OI����DF�_L�0�r�Q�PLM��F^�HRDYO,�af�RG��H���a�|0p�/�MULSE������Qp�$J�xzJ�r�w�{FAN�_ALMp���WR=N��HARD�0�VZ0P]R�2���A���e_��fAU�R�ȴRTO_SBR &E�O`#��ӓ��;�_MPINFQ���N��Y�REG�6NQV�Pf3�fDA@N��sFL����$M�� ��`S����P�����CMѐNF-��1����h��A��0$Δ1$Y oQ�b�Q�0�� ���cEG�0+c`p+A1R=`CHu25Rr:�T��eAXEEgRO�BBjREDBfWRd,� q_�$sSY�`�ep�S�WRI,�>�STr@CcP�p�pE��0G6�Rr��;`B� R��7\��2�OTOi��0��ARYBc4~�2�̹"t`FI�`�c$�LINK�GTH�S�PT_�R�rF8Rr|XYZ�R:�9�OFFZ�S){o8B@`����/��@�P�FI@1�����CXt��Zd_J�A�R�r`����30Rr�@�*!dm�b"CFA�eDUn�rHu3����TUR��!X�ӛ%BI�X� `�J'FL|�a�8 � ԝ�	3ʡg� +1��0Kg`M�d�&�Qs�����°�pSOR�Q&�Oa�P(���`O � �1ɐj4��Ma��~4'OVE�1MIPk1 ��5�5�6_Q�70c��7��4ANڡV �1���1�`�0�k1 �5�1�7(E(E�3OaSERla�	��E,�H�P��fDAA�P����!�@o�l�o�AX /��Ro�2��U�EQ� �I{��I���JN �J��J$�J��J��J1 [ �F/��I/��I/��I /��I/�Y/�Y/�(Y�/�8Y/�HYeQYYDEBUڣ$����I�	ao�wABo�m��qr3Vb�٢ 
$b �LeʡXgQqXg�� XgNXgXg$Xg��Xg���g ��U�L�AB�J5֠�G�RO[�J"��K�B_/�MF��s� �v�5qK51u�=vAND 0��[DL��^A�zw K���� �x1ѝxN��NT��#��pVEL5��4�qm��x9���NA��V�$���ASS  �����* *  ��_�SI@���#��)�I�Y�n��(�AAVM���K 2 T�� 0 � �5�����\���� ��	݀΍�* U��ߏ��!�͌@�L�܁R��������e�BS�1  �16�� <u����
��.� @�R�d�v��������� Я�����*�<�N� `�r���������̿޿ ���&�8�J�\�n� �ϒϤ϶��������� �"�4�F�X�j�|ߎ� �߲��������߱��p�MAX/� ����ʓ  d�IN��*��PRE_EXE;�g�J�!43���T�e�IOCNV,�"<� �&�P��a �;�Ɨ��IO_�� �1r�P $b��`���V���U�?��� ��$�6�H�Z�l�~� ��������������  2DVhz�� �����
. @Rdv���� ���//*/</N/ `/r/�/�/�/�/�/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�?�? O"O4OFOXOjO|O�O �O�O�O�O�O�O__ 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o Poboto�o�o�o�o�o �o�o(:L^ p�������  ��$�6�H�Z�l�~� ������Ə؏����  �2�D�V�h�z��������ԟ����LA�RMRECOV �~�!�J���LM_DG ����� �LM_IF ��+��ߥ���ɯۯ�骓���0�B�S�, 
 S�|���@�����ƿؿ�$�� ���1��U�g�yϋ�����NGTOL � ~� 	 A�   �����PPINFO Z� Y��*�<�N�!�  f�P�~�?�m� �ߑ��ߵ������%��5�[����χ�� �����������)��;�M�_�m�PPLI�CATION ?}���H��Handl�ingTool ��� 
V9.1�0P/30��j�?
88340�����F0����1028��������7DF�1��j���None�j�FRAj� �6w�_ACoTIVE�  �����  �UTOMOD� ^��Ê�CHGAPONL�� �OUPL�ED 1��� �
 2�CU�REQ 1	�� � T<<<	�����@��<�����Hk�HTTHKY�A�o�� �////�/S/e/w/ �/�/�/�/�/�/�/? ?+?�?O?a?s?�?�? �?�?�?�?�?OO'O �OKO]OoO�O�O�O�O �O�O�O�O_#_}_G_ Y_k_�_�_�_�_�_�_ �_�_ooyoCoUogo �o�o�o�o�o�o�o�o 	u?Qc�� �������� q�;�M�_�}������� ��ˏݏ���m�7� I�[�y��������ǟ ٟ����i�3�E�W� u�{�������ïկ� ���e�/�A�S�q�w���NTO����DO_CLEAN�|��NM  �� <_�qσϕ����BDSPDRY�RϊHI� ;�@ L��%�7�I�[�m�߀�ߣߵ������߇MAX~�������	��X���PL�UGG� ���P�RC��B9�=�����c�Oh�����SEGF� K������ 9�K��%�7�I�[�����LAP������ ��������	-?�Qcu��TOT�AL+�T��USE+NU��� ޸���NRGDISPWMMC��0�C��&�@@���O�������_STRI�NG 1
�
��M� S�
�
^_ITEM1h  n���� ����//&/8/ J/\/n/�/�/�/�/�/��/I/O S�IGNALb�Tryout M�odeiInp�0Simulat{edmOut,<OVERR��� = 100lIn cycl 5�mProg A�bor63m4S�tatusk	H�eartbeat�gMH Fauyl�7�3Aler�9 �/�?�?�?O#O5OGO8YOkO}O ��d ��v�O�O�O�O__ (_:_L_^_p_�_�_�_��_�_�_�_ oo�OWOR��dJa�O$oro �o�o�o�o�o�o�o &8J\n��8���~POb�1 �pbk��#�5�G�Y� k�}�������ŏ׏� ����1�C�U�g��rDEV�~������ ˟ݟ���%�7�I� [�m��������ǯٯ�����PALT �M6�bo�^�p����� ����ʿܿ� ��$� 6�H�Z�l�~ϐϢ�$�GRI�d��N��� ��&�8�J�\�n߀� �ߤ߶���������� "�4�F���� R�M~� ��X��������� � �$�6�H�Z�l�~��������������l�PREG:�# ����J\ n������� �"4FXj|���-�$ARG_�J`D ?	������ � 	$�&	+[�]���')��SBN_CONGFIG� �$1#2�=!!CII_S?AVE  �$F!�9#�TCELLSETUP ��%  OME_I�O�-�,%MOV�_H� �/�/REP����/�UTOBA�CKv!�@"�FRA:\ ��/F '`�0�C8� T;? � 23/0�7/18 17:_50:04(��?�?�?�?4<�� O6OHOZOlO~O�O�$O�O�O�O�O__ �O<_N_`_r_�_�_�_ 3_�_�_�_oo&o�_ Jo\ono�o�o�o�o��ׁ  /1_3_\�ATBCKCTL.TM���o+\=;INI9�v5�6%J!0MESSA�GV dqF!�o{ODGE_D� Y&6%�x�O���3PAUS�� !�� , 	� ���,		�8�"� \�F�X���|����� �֏����F��t�p?TSK  �}C?<I0UPDT�pbw�d���vXWZD�_ENBbt2*��S�TAau����XI�S$ UNT 2��C!E � 	 �8�� ������!D � �p� �/"
T���.�������
9�r���F������/6�5��5 [^. 8��a�¯����\����MET��2i��b# P�B���A�-mA�J� 7MWAA%���A��٭>a�:>ٻ�>p��35ؔ>B��>H�0�S�CRDCFG 1��%1 �^%C"篻�Ϳ߿���<?
QZ)��e� wωϛϭϿ�&���J� ��+�=�O�a�����1GR��������`NA� �	�4��_ED`p1z���_��%-�`EDT-���*�B�Y�b?$� -3�
�"O�&
��  ����2��#� �G��_���G����6����3��+]��� ̔\��Z�l�����4K�������t@�&8�\��5 �d���@���(��6�S0/w ��/w/��f/���7�//�/C/���/C? �/�/2?�/��8{?���?�f&��?OV?h?�?�?��9GO�?�O�?i&�pO�O"O4O�OXO��CR���/__q_ = :_�_�O�O�_"_����?NO_DEL�ߞ��GE_UNUSE��ߜ�IGALLO�W 1��  � (*SYS�TEM*֣	$SERV_GR�k�_`�pREGhe$8�c֬_`NUM�j�c��mPMU`֥�LAY�֬?PMPALap�e�CYC1p��c }x�`�n%sULSU�o0�mr�qjcL;tt�BOXORI�eC�UR_ap�mPM�CNV�fap1�0~�pT4DLI�ǐZ|i	*PRO�GRAgdPG�_MI�n�)�AL(�u6� �)�BT�_n�$FLUI_RESUw���o��Ä#MRvn�`�\�_Β ��+�=�O�a�s��� ������͟ߟ��� '�9�K�]�o������� ��ɯۯ����#��R�LAL_OUT �Nk���WD_�ABORp/o��I�TR_RTN  ��D��ل�NONgSTO�Я� 8h�CE_RIA_IL,`�������FCFG ��x�ĨN�_LIMvb�2�� �  �� 	��gϳB<�҄��e�@�  VϷ����ϨH
�����2�PAn�GP ;1�ޥ��n߀ߒ�Q�C>  )C.���f��z���ߪ�Ї�Б�Ж�Р
�Ъ�д�Թ������������C���ǀW CѶ��J��G�?��HE�PON�FIπ��d�G_Pv�p1;� �U ;ծ�����������|,�d�KPAUS~q31;��� �r.� t�;�b����������� ����0@fL�����6�M��N�FO 1?�� �T��B��̵��5�Au�9	�]��Ǝ�@���K D5Oy����C����($6�T5�+��P� �8�h�Ca����.~:��1ﯼ���O��ϨG��COLL/ECT_�?�x�ǯEN�p�����n�NDE�?��;c�R1234?567890'�B ya�//&��HC��C)j/�/y\i/{/�/z[ �/�/?�/�/?`?+? =?O?�?s?�?�?�?�? �?�?8OOO'O�OKO ]OoO�O�O�O�O_�Ot�9�� �>�IO !)������_�_�_�_`W[TR6�2"D](�b{Y
�O�^o�#o]x jt�i_MOR9��$;� ��:B��\`�e �i�o�o��o�o�o�kbb1�:�%
pm,t�?]�]���>qR�KFt�`�R��&�utqtrC4 W A�����x�SA����B�pCd �B��d C  @�r��q�:d�TQbZqI#'d}?�s�9�(pm����dZqTo_DEFB� {�%oR��thPNUS�E��s���g�KEY?_TBL  �������	
��� !"#$%&�'()*+,-.�/(':;<=>?�@ABC)�GHI�JKLMNOPQ�RSTUVWXY�Z[\]^_`a�bcdefghi�jklmnopq�rstuvwxy�z{|}~����������������������������������������������������������������������������,���͓���������������������������������耇�������������������s��4Q��LCKp�8ٹ��p�STA���t�_AUTO_DOrζkv�IND�<ٞ�R_T1��旃T23�ݵʳ��T{RL(�LETE���z�_SCREE�N ;�k�csc�UʰMM�ENU 1)l� <7�@������ F��#�I���Y�k��� �����ſ׿��6�� �l�C�UϢ�yϋϱ� ������ ���	�V�-� ?�eߞ�u߇��߽߫� 
������R�)�;�� _�q��������� ��<��%�r�I�[��� ������������&�� 5nEW�{� ����"�X /A�ew����/)\ʠ_MANgUALo�*�DB'a�.b����DBG_E7RRL.�*֫�Q� /�/�/�.~L!NUMLIM����lu
L!PXW�ORK 1+֫��/#?5?G?Y?k?mD�BTB_�� ,�{-�s�Qst3QD�B_AWAYT#ޅQGCP lr=�9��"�2_AL� ٟ��2P"Yn���lpE(_�n  1-�[,p
�?POJf@O}O�6_M&�IS֐�;@�p�C�ONTIM���&lt��FI
� CMOTNENDt��DRECORD ;13֫ ��OxsG�O�KQ9_x{�2 w_�_�_�_DX�_�_K_  oo_$o6oHo�_�_~o �_�oo�o�o�o�o�o  �oD�ohz�� �1�U
��.� @��d��������� Џ�Q��u����N� `�r���󏨟���;� ���&���J�5�C� �����ȯ7��ׯ m�"���F�X�j��y� ���Ŀ3����ϣ� ��Bϱ�f�տ�ϜϮ� ��[���S��w�,�>��P�b��Ͽ2TOLEoRENC�4B�B��0L��L CSS�_CNSTCY +249�Y e�B����������#�5� G�]�k�}�����������������DEVICE 25�� �6o������� ��������&�O���HNDGD 6�۬0Cz9
Q��_LS 27Y�8 �����:���PARAM �8,I�2�5&�ySLAVE 9Y�E_CFG :�F&dMC:�\��L%04d.'CSV%@c�B6�A �CH kAkO&/B/X�&�2"_!o/])\!1@�JPя#N.A�1�n_CRC_OU�T ;Y��1*__NOCODz<,G��SGN =�"UR#M��20-JUL-23 02:57��0A18>517�:51�~� V�hr9n1&o0�61�M��Þ��j��1�>�V�ERSION �):V4.2�.11�KEFLO�GIC 1>�� 	�(1@I�!�M�2PROG_E�NB Xa=CULS��G `�2_AC�CLIM�F����|CWRST�JNT�G
S���1M�OFLX!2�DINI�T ?��"U�� ��FOPTu ?�	�F�B
 	�R575&'P74j,Y6-X7-W50QX�4WR2-T�({_�7
TTO  ]�?�_��6V�@DEX�Gd��B� �SPATHw A):A\�_�5oGo|�HCP_CLNTID ?�6� �+Ӈo���IAG_GRP� 2D� �� 	 D��  D�� D�  B��Т��ff�j�`���o�l�a��%��B��N�C�-B�z��Bp��e�`�imp2m�7 789012�3456xq�G�`��  Ao�
�Aj{Ad�]�AW�AP���AJ=qAC�33A<�4zᘝj�p�!@��]pA,�q��A�����B4�lf�dX�!�
�ru�ppQ�A�j�HAeG�A}_�pY��AS�p�M2�F�RA@(��J���t�J��I��@�p������?��@��HL�^�pp��������33<���=q@~�R@�xQ�@q�@�k�@dz�@]��Vff؏����� ���s>�l�Ϳ@e@^J�W�
=@Pv�G��@@v�7ڐ.{@d�v���������S>��M���AR�<(��@5Ґ/\)@(/��@!R�֏ � �$�6��ĭ���ܯ "�4����V�|�Z��� ��<�N�������0� B�̿R��B�`�r5����M�ّe��m>��R>��?�33?9�������m7'Ŭz��6��4�F��7��L�m@ž����ڐ␀N�Њ=�@�pAh������c= c<���]>*�H>�V>�3�>�����m<���<�b�a�i�L. �?�� �C�  <w(�UX" 4��A�>��ё��ٝiA�� ?�el���t���� ,��H��8�b���r���z����x�?�7���>�(�>!ʽ���=����m�7�G��G��m�����I��m����i�@��Ҁ�@Q�?L��Ly�o�g�v\��
��]p'�@����8����	�gC� ���Cu��Zl� <� ���`���&%�18�� ����4�J6�<�D�5OL��rC��� �5�qW�(S���$�z��	�($6�T��Á�i���x������{�ʝm;��t���9/�aCT_CONFIG E?>i3eg�%�a�STBF_TTS�G
UI�#�0�C�A�&� MAU�@JOJ"�MSW_CFX F�k  �p�:OCV7IEW� G�-�a���o=?O?a?s?�? �?�B+?�?�?�?�?O O�?>OPObOtO�O�O 'O�O�O�O�O__(_ �OL_^_p_�_�_�_5_ �_�_�_ oo$o�_Ho Zolo~o�o�o�oCo�o �o�o 2�oVh`z���@,RC�#{��"!L�~����A�0�e�T����$SB�L_FAULT �I�z 8��GPM�SK�'��L TDI�AG J\)�!���1�UD�1: 6789012345�p"1�j'�uP&/O�a�s��� ������͟ߟ��� '�9�K�]�o�����y���
>���F&TRECP���
���%� ��=�:�L�^�p����� ����ʿܿ� ��$� 6�H�Zρ�������7�UMP_OPTIcON� ����TR�"t�#����PME�%���Y_TEMP � È�3B�̞ 1��A.��UN�I� �%1��&YN_?BRK K?6?EDITOR�����
��_ԠENT �1L�y  ,�&PART1 TLOG ����f����2���&M�AI���߫�&OMAY��[���F� �߇���� u���J������
IRVWA�I����&-BC?KEDT- ��/����PICKSIM_��[���y���o"�x����������� ��3WiP� t�������~�MGDI_STaAD� !1�y�NC7;1M�+ �`�r��
��d���� �/!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?��j?|?�? �?�9��?�?�?�?
O O.O@OROdOvO�O�O �O�O�O�O�O__*_ <_�:c?m__�_�_�? �_�_�_�_o!o3oEo Woio{o�o�o�o�o�o �o�o/A[_e w���_���� ��+�=�O�a�s��� ������͏ߏ��� '�9�SA�o������ ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�K�]� g�y���A�����ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�C�U�_�q߃ߕ� ������������%� 7�I�[�m����� ���������!�3�M� W�i�{����߱����� ����/ASe w������� +E�Oas� �������// '/9/K/]/o/�/�/�/ �/�/�/�/�/?#?= /?Y?k?}?���?�? �?�?�?OO1OCOUO gOyO�O�O�O�O�O�O �O	__5?G?Q_c_u_ �_�?�_�_�_�_�_o o)o;oMo_oqo�o�o �o�o�o�o�o�_ ?_I[m�_�� �����!�3�E� W�i�{�������ÏՏ �����7A�S�e� w��������џ��� ��+�=�O�a�s��� ������ͯ߯��� /��K�]�o������ ��ɿۿ����#�5� G�Y�k�}Ϗϡϳ��� �������'�9�C�U� g�ߓ��߯������� ��	��-�?�Q�c�u� ������������ �1�;�M�_�q��ߕ� ����������% 7I[m��� ����)�3E Wi������� ��////A/S/e/ w/�/�/�/�/�/�/�/ ?!+?=?O?a?{m? �?�?�?�?�?�?OO 'O9OKO]OoO�O�O�O �O�O�O�O�O?_5_ G_Y_s?�?�_�_�_�_ �_�_�_oo1oCoUo goyo�o�o�o�o�o�o �o_#_-?Qc}_ �������� �)�;�M�_�q����� ����ˏݏ�i%� 7�I�[�u������� ǟٟ����!�3�E� W�i�{�������ïկ �����/�A�S�m� w���������ѿ��� ��+�=�O�a�sυ� �ϩϻ���������� '�9�K�e�[߁ߓߥ� �����������#�5� G�Y�k�}������ �������1�C��� o�y������������� ��	-?Qcu ��������� );Mg�q�� �����//%/ 7/I/[/m//�/�/�/ �/�/�/?!?3?E? _i?{?�?�?�?�?�? �?�?OO/OAOSOeO wO�O�O�O�O�O�O�/ __+_=_W?I_s_�_ �_�_�_�_�_�_oo 'o9oKo]ooo�o�o�o �o�o�o�O�o#5 O_a_k}���� �����1�C�U� g�y���������ӏ�o �o	��-�?�Yc�u� ��������ϟ��� �)�;�M�_�q����� ����˯E�����%� 7�Q�[�m�������� ǿٿ����!�3�E� W�i�{ύϟϱ����� �����/�I�S�e� w߉ߛ߭߿������� ��+�=�O�a�s�� ������������ '�A�7�]�o������� ����������#5 GYk}������� �$ENETMODE 1NB���  �������� RROR_PR_OG %�
%���an<TABLE  �L������<SEV_N�UM 
  �� <_A�UTO_ENB � (9_NON! O� "_  *�Y �Y %�Y �Y  +X r/x�/�/2$FLTR/0&HIS���++_ALM 1P�� ���Y,��+�/2?D?V?h?z?�?r�/_�8   ��W!�:� TCP_VER !�
�!Y�?$EXTL�OG_REQ�&9�))#CSIZ,OD�STKIIG%�~ BTOL  ��{Dz�"�A D_BWD�0�@�&�A�#�CDI�A QB��C��KSTEP�O�O� �@�OP_DOkO�F�ACTORY_T�UN�'d3YDR_?GRP 1R�	�!�d 	�?�_{P��*u����RHB ��2 ���� �e9 ����V{S�_�]{P�B���B�F>�C��B���AԂ=Bu� ��[A���B��B��A����AI��B ��]�_WoBo{ofo�o��o�o�o  @��:A|=@9q���o��
 F��5W&b�`��A�$ � #�4<�o`K�n�Y�  �qA��`w�33�r�33�]/@UUT�z@�`�p�j$>u.�>*���<����]E�� F@ ��p&��]J��NJ�k�I'PKH�u��IP�sF�!���]?�  �j��9�<9��896C�'6<,5����~����=����a��� �_&���#�tFEATURE� SB��@"�HandlingTool 	����Engli�sh Dicti�onary�4Dw St��ard	���Analog �I/O@�I�gle� Shift\�u�to Softw�are Upda�te��matic Backup����ground �Edit��Ca�meraW�F[�CnrRndIm����ommon calib UI���n͑�Moni�tor&�tr�R�eliabp��D�HCP�]�ata Acquis5�~^�iagnos���T�x�ocument VieweA��`�ual Che�ck Safet�y!��hance�d!����sʠFr�ސ�xt. DI�O 1�fi��&�e�nd��Err@�L(��B��sA�rR�1�� �@�FCTN /Menu�v\����TP In��fayc���GigE���εƐp Mask� Exc��g#�H�T��Proxy �Svˤ�igh-wSpe��Ski��Ŧ�5�mmuni�c��ons<�urࡰ��s�X���con�nect 2s�n{cr��stru#�$qʚ�e��۠J����KAREL Cmod. L �ua�~��Run-Ti"��Env�Ȅ�el u+��s��S/W�Licenseݣ�ʬX�Book(S�ystem)�M�ACROs,3�/�Offsew�V�H05���q�[�MR:�6����MechStoEp�t����V�iS��s���x��T�����o}dq�witch���ӡ�.{��Optqm,���filʬ��gi�V�ulti�-T��Г�PCMO fun�Ǣ�o��xޢ����RegiK�YrW���riàF�����U�Num Se�l��� � Adj�uG��=�s�N�ta�tu��f�Ū�RDM Robot ��scove)���e�a��"�Freq �AnlyW�Remļ�5�n7�����Se�rvo5���SN�PX b�x�SN���Cli¡%t�LGibr(�E�� ���W o0�t��ss#ag����0 ��n����0/I���MI�LIB��P F�irm���P��A�ccǐϛTPTXm��elnn���x�jղorquq�imula?��bu�PaѱƐZ�:(�&�ev.����ri۠:USB� port �i�PL�aà�R E�VNT��nexcept�������,��VC�rR�I���V��o"�%Wz+�S8 SC4�/SG�E�/�%UI�Web Pl}� >i��'4�����x�ZDT ApplP��&�?|7Grid��p�layv=� ���7R�f".7��6���/Y�-10iA/8L�?�Alarm C�ause/��ed>*�Ascii�<��Loadʠ:JUp�lP@�l�7�Gu�=�rO�BP��Ֆyc�p�����蠕�RAp� �9�NRTJ��On�e Hel��漿������1�tr;�ROS E�th
�t�BeW7i}R�$2D Pk;�uVIm+�Fd�� �^�nsp���Q�64MB DRAM�O��SFRO�_ېellW��shao g�cK�e��p�2ltyp�s'�ԗ�B��D�.�maiܠ;�(��T�qV�R7��FL!PSup�c���8 pL���cro~����W�4��&��auestz&rtڡ���/�3DL}|�Q���T�y,K��l Buiz��n�/APLC�2�uVZ��/CGl��'CRG#��$D��@�fR�LS[��%BUw�b�%Kі��!TA����B�,يE�TCB��ʏ��/��^�TC��v��%��TEHǟٖ"�ؗ!V�����/��F�H����G:���n�����2��H¯��IA߯�Lޯ��LN���M�� D���D�����N���!P��������RR���!Sڿ�����W.�@ǜ���$VGFf�x�P�2Z���2��ǂϔ�B$�ϔ�D�ϔ�Fr������"TUT��01�J�\�2f�\�TBGyG��rain��sUI*ЦUHMI��r ponU2�8���a�f{ �R�v�VKAR3EL��_TP� ��e��R9�0�B�o�f� x������������ �5�,�>�k�b�t��� ������������1 (:g^p��� ���� -$6 cZl����� ���)/ /2/_/V/ h/�/�/�/�/�/�/�/ �/%??.?[?R?d?�? �?�?�?�?�?�?�?!O O*OWONO`O�O�O�O �O�O�O�O�O__&_ S_J_\_�_�_�_�_�_ �_�_�_oo"oOoFo Xo�o|o�o�o�o�o�o �oKBT� x������� ��G�>�P�}�t��� ����׏Ώ����� C�:�L�y�p������� ӟʟܟ	� ��?�6� H�u�l�~�����ϯƯ د����;�2�D�q� h�z�����˿¿Կ� ��
�7�.�@�m�d�v� �Ϛ��Ͼ�������� 3�*�<�i�`�r߄ߖ� �ߺ��������/�&� 8�e�\�n����� ��������+�"�4�a� X�j�|����������� ����'0]Tf x������� #,YPbt� ������// (/U/L/^/p/�/�/�/ �/�/�/�/??$?Q? H?Z?l?~?�?�?�?�? �?�?OO OMODOVO hOzO�O�O�O�O�O�O _
__I_@_R_d_v_ �_�_�_�_�_�_oo oEo<oNo`oro�o�o �o�o�o�oA 8J\n���� �����=�4�F� X�j�������͏ď֏ ����9�0�B�T�f� ������ɟ��ҟ���� �5�,�>�P�b����� ��ů��ί����1� (�:�L�^��������� ��ʿ��� �-�$�6� H�Zχ�~ϐϽϴ��� ������)� �2�D�V� ��zߌ߹߰������� ��%��.�@�R��v� �����������!� �*�<�N�{�r����� ����������& 8Jwn�������  �H552��21nR7850�J614ATU]P)545)6�VCAMCRIndUIF)28e�NRE52XR�63SCHDwOCV�CSU�869)04EI�OC�4R69�XESETAWJ�7WR68MA{SKPRXY}]7OCO(3Ah! (3`&J6'�53�H�(LCH^H&OPLGA0x&�MHCRI&S�'MkCS@0$'554�MDSW!7k'OP�k'MPRl&��(0n(PCM|R0g7�! 4� �'51L5u1�80LPRS'�69`&FRDdFwREQMCN{93(SNBA�^�'SHLBFM'Gt�82(HTC@�TMIL�TP�A�TPTXYFEL�6� �8wJ95�TUTl'�95`&UEV&U�ECH&UFRdV�CC XO�&VIP�dFCSC�FCSGt��IWEB@7HTT@R6��H�CG_WIGGWIP�GS�VRCdFDGvk'H7�R66L�R7'R�8R53V�768�82x&R�*�4�W664R64nNVD&R6�'`9 �X�9 �D0+g�F~hCLIP8KC�MS��`@STY�$WTO@NN`&OkRS�&M�8OL�hWENDLWS�hwFVR�V3D$X�{PBV�FAPL��APVl&CCGn@CCR�&CDWwCDL�VCSB��CSK,6CT{GC#TBHV�p�hC(F�p�xC<WTC|�ppw�TC�wTC&CT1E�9�|wTE�9�V0WTF�xF�hG�x)Gx�$�H$�IF��\$��GCTM�hM�UM�xN$�P��P�xYR�x�hTS�xW8�n�VVGFP�P2 W�P2�6e�\�B\�D�\�F|VP��VT���VTB�wV��IHWGV�P՗K$WV_V��)�;�M� _�q���������˯ݯ ���%�7�I�[�m� �������ǿٿ��� �!�3�E�W�i�{ύ� �ϱ����������� /�A�S�e�w߉ߛ߭� ����������+�=� O�a�s������� ������'�9�K�]� o��������������� ��#5GYk} ������� 1CUgy�� �����	//-/ ?/Q/c/u/�/�/�/�/ �/�/�/??)?;?M? _?q?�?�?�?�?�?�? �?OO%O7OIO[OmO O�O�O�O�O�O�O�O _!_3_E_W_i_{_�_ �_�_�_�_�_�_oo /oAoSoeowo�o�o�o �o�o�o�o+= Oas����� ����'�9�K�]� o���������ɏۏ��  H5�5Ȕ�����R7�8�50	�J61�4	�ATU�?�5�459�6	�VCA�M	�CRI��UI�F9�28��NREv�52x�R63��SCH	�DOCV���CSU�869z9�0H�EIOCɛ�4(�R69x�ES�ETY�w�J7w�R{68�MASK	��PRXY��7	�OCOy�3Y�(���8�m3تJ67�53(��H�LCH��OP�LGY�0��MHCuR��Sw�MCSX��0��55H�MDS�Wٻ�OP�MP�R��(�08�PCM��R07˅�H����(�51h�51x�0nh�PRSx�69ت�FRD��FREQn�MCN	�938��SNBAٛ�SH�LB	�M7��ȼ2�8�HTCX�TMI�L�(�TPAH�T7PTXy�EL�ʅ��(�8'�%��J95n��TUT�95تwUEVx�UEC��wUFR��VCCX��O��VIP��CS�C��CSGȚ�I�	�WEBX�HTTfX�R6ל��CG��{IG��IPGS	��RC��DG�H7n'�R66h�R7g��Rv�R53h�68�h�2��R6�4��6�6H�R64�NVDx�R6����h��������D0��FVCsLI�g�CMSH�ܕ X�STY��TOvX�NNتORS���M��OL�END��Lg�S�FVR�H�V3D�짛PB�V��APLH�AP�V�CCGX�CC�Rx�CDg�CDL�(�CSB�CSKv�CT��CTB��D �C8�5 ,C��cTC��5 �TC�;TCx�CTE��� ƨTE�� ��TF*,F�G,G�-�,�H�,I�E0�,��C�TM�Mx,M�N*�,PH<P,R,��TS,W�=(�VGmFKP2X�P2��T5@(LB(LD(LF��VPW;VT��@(��VTB�V�IHRw�V5��KK��V�� �_1_C_U_g_y_�_ �_�_�_�_�_�_	oo -o?oQocouo�o�o�o �o�o�o�o); M_q����� ����%�7�I�[� m��������Ǐُ� ���!�3�E�W�i�{� ������ß՟���� �/�A�S�e�w����� ����ѯ�����+� =�O�a�s��������� Ϳ߿���'�9�K� ]�oρϓϥϷ����� �����#�5�G�Y�k� }ߏߡ߳��������� ��1�C�U�g�y�� �����������	�� -�?�Q�c�u������� ��������); M_q����� ��%7I[ m������ �/!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?e?w?�?�? �?�?�?�?�?OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_K_ ]_o_�_�_�_�_�_�_ �_�_o#o5oGoYoko }o�o�o�o�o�o�o�o 1CUgy� ������	�� -�?�Q�c�u�������轏Ϗ��S�TD�LANG�� �2�D�V�h� z�������ԟ��� 
��.�@�R�d�v��� ������Я����� *�<�N�`�r������� ��̿޿���&�8� J�\�nπϒϤ϶��� �������"�4�F�X��j�|ߎߠ߲�RBT�OPTN�����߀���#�5�G�Y�k�DPN�������� ������%�7�I�[� m�������������� ��!3EWi{ ������� /ASew�� �����*�/ 1/C/U/g/y/�/�/�/ �/�/�/�/	??-??? Q?c?u?�?�?�?�?�? �?�?OO)O;OMO_O qO�O�O�O�O�O�O�O __%_7_I_[_m__ �_�_�_�_�_�_�_o !o3oEoWoio{o�o�o �o�o�o�o�o/ ASew���� �����+�=�O� a�s���������͏ߏ ���'�9�K�]�o� ��������ɟ۟��� �#�5�G�Y�k�}��� ����ůׯ����� 1�C�U�g�y������� ��ӿ���	��-�?� Q�c�uχϙϫϽ��� ������)�;�M�_� q߃ߕߧ߹������� ��%�7�I�[�m�� ������������� !�3�E�W�i�{����� ����������/ASe�h�������99���$FEAT_AD�D ?	����  	�%7I[m �������/ !/3/E/W/i/{/�/�/ �/�/�/�/�/??/? A?S?e?w?�?�?�?�? �?�?�?OO+O=OOO aOsO�O�O�O�O�O�O �O__'_9_K_]_o_ �_�_�_�_�_�_�_�_ o#o5oGoYoko}o�o �o�o�o�o�o�o 1CUgy��� ����	��-�?� Q�c�u���������Ϗ ����)�;�M�_� q���������˟ݟ� ��%�7�I�[�m�� ������ǯٯ���� !�3�E�W�i�{����� ��ÿտ�����/� A�S�e�wωϛϭϿ���������DEM�O S   �N�D�V߃� zߌ߹߰��������� ��I�@�R��v�� ������������ E�<�N�{�r������� ��������
A8 Jwn����� ��=4Fs j|������ //9/0/B/o/f/x/ �/�/�/�/�/�/�/? 5?,?>?k?b?t?�?�? �?�?�?�?�?O1O(O :OgO^OpO�O�O�O�O �O�O�O _-_$_6_c_ Z_l_�_�_�_�_�_�_ �_�_)o o2o_oVoho �o�o�o�o�o�o�o�o %.[Rd�� ������!�� *�W�N�`�������Ï ��̏�����&�S� J�\�����������ȟ ����"�O�F�X� ��|�������įޯ� ���K�B�T���x� ��������ڿ��� �G�>�P�}�tφϳ� �ϼ��������C� :�L�y�p߂߯ߦ߸� ����	� ��?�6�H� u�l�~�������� ����;�2�D�q�h� z������������� 
7.@mdv� ������3 *<i`r��� ����///&/8/ e/\/n/�/�/�/�/�/ �/�/�/+?"?4?a?X? j?�?�?�?�?�?�?�? �?'OO0O]OTOfO�O �O�O�O�O�O�O�O#_ _,_Y_P_b_�_�_�_ �_�_�_�_�_oo(o UoLo^o�o�o�o�o�o �o�o�o$QH Z�~����� ��� �M�D�V��� z�������ݏԏ�� 
��I�@�R��v��� ����ٟП���� E�<�N�{�r������� կ̯ޯ���A�8� J�w�n�������ѿȿ ڿ����=�4�F�s� j�|ϖϠ�������� ���9�0�B�o�f�x� �ߜ������������ 5�,�>�k�b�t��� ����������1�(� :�g�^�p��������� ������ -$6c Zl������ ��) 2_Vh �������� %//./[/R/d/~/�/ �/�/�/�/�/�/!?? *?W?N?`?z?�?�?�? �?�?�?�?OO&OSO JO\OvO�O�O�O�O�O �O�O__"_O_F_X_ r_|_�_�_�_�_�_�_ oooKoBoTonoxo �o�o�o�o�o�o G>Pjt�� �������C� :�L�f�p�������ӏ ʏ܏	� ��?�6�H� b�l�������ϟƟ؟ ����;�2�D�^�h� ������˯¯ԯ��� 
�7�.�@�Z�d����� ��ǿ��п�����3� *�<�V�`ύτϖ��� ���������/�&�8� R�\߉߀ߒ߿߶��� ������+�"�4�N�X� ��|���������� ��'��0�J�T���x� ��������������# ,FP}t�� �����( BLyp���� ���//$/>/H/ u/l/~/�/�/�/�/�/ �/?? ?:?D?q?h? z?�?�?�?�?�?�?O 
OO6O@OmOdOvO�O �O�O�O�O�O__2]  )XH_Z_ l_~_�_�_�_�_�_�_ �_o o2oDoVohozo �o�o�o�o�o�o�o
 .@Rdv�� �������*� <�N�`�r��������� ̏ޏ����&�8�J� \�n���������ȟڟ ����"�4�F�X�j� |�������į֯��� ��0�B�T�f�x��� ������ҿ����� ,�>�P�b�tφϘϪ� ����������(�:� L�^�p߂ߔߦ߸��� ���� ��$�6�H�Z� l�~���������� ��� �2�D�V�h�z� ��������������
 .@Rdv�� �����* <N`r���� ���//&/8/J/ \/n/�/�/�/�/�/�/ �/�/?"?4?F?X?j? |?�?�?�?�?�?�?�? OO0OBOTOfOxO�O �O�O�O�O�O�O__ ,_>_P_b_t_�_�_�_ �_�_�_�_oo(o:o Lo^opo�o�o�o�o�o �o�o $6HZ l~������ �� �2�D�V�h�z� ������ԏ���
� �.�@�R�d�v����� ����П�����*� <�N�`�r��������� ̯ޯ���&�8�J� \�n���������ȿڿ ����"�4�F�X�j� |ώϠϲ������������0�   1�6�L�^�p߂ߔߦ� �������� ��$�6� H�Z�l�~������ ������� �2�D�V� h�z������������� ��
.@Rdv ������� *<N`r�� �����//&/ 8/J/\/n/�/�/�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�o�o $6 HZl~���� ���� �2�D�V� h�z�������ԏ� ��
��.�@�R�d�v� ��������П���� �*�<�N�`�r����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ����� ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������ (�:�L�^�p������� �������� $6 HZl~���� ��� 2DV hz������ �
//./@/R/d/v/ �/�/�/�/�/�/�/? ?*?<?N?`?r?�?�? �?�?�?�?�?OO&O 8OJO\OnO�O�O�O�O �O�O�O�O_"_4_F_ X_j_|_�_�_�_�_�_ �_�_oo0oBoTofo xo�o�o�o�o�o�o�o ,>Pbt� �������� (�:�L�^�p������� ��ʏ܏� ��$�6� H�Z�l�~�������Ɵ ؟���� �2�D�V� h�z�������¯ԯ� ��
��.�@�R�d�v� ��������п���� �*�<�N�`�rτϖ� �Ϻ���������&�
5�:�-�P�b�t� �ߘߪ߼�������� �(�:�L�^�p��� ��������� ��$� 6�H�Z�l�~������� �������� 2D Vhz����� ��
.@Rd v������� //*/</N/`/r/�/ �/�/�/�/�/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FOXOjO|O�O�O�O�O �O�O�O__0_B_T_ f_x_�_�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o (:L^p�� ����� ��$� 6�H�Z�l�~������� Ə؏���� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4� F�X�j�|ߎߠ߲��� ��������0�B�T� f�x���������� ����,�>�P�b�t� �������������� (:L^p�� ����� $ 6HZl~��� ����/ /2/D/ V/h/z/�/�/�/�/�/ �/�/
??.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O�O�O�O�O�O__�&_8Y�$FEAT�_DEMOIN [ =T�hP�=P}PTINDEX][�lQ�PPILEC�OMP T�;���QkRKU��PSETUP2 �U�U�R��  N �Q�S_A�P2BCK 1V~�Y  �)9XDok%�_:o=P�P (oeo;U�_�o o�oDo �o�ozo�o3E�o i�o��.�R� ����A��N�w� ���*���я`����� �+���O�ޏs���� ��8�͟\�ڟ���'� ��K�]�쟁������ F�ۯj������5�į Y��f������B�׿ �x�Ϝ�1�C�ҿg� ���ϝ�,���P���t� ��ߪ�?���c�u�� ��(߽���^��߂�� )��M���q� �~�� 6���Z������%��� I�[���������D� ��h�����
3�Y�P�P�_ 2�P*�.VR:���*��������n P�C���FR6�:�4�X�T |P|�y�_PI<���*.Fq/"��	�<,�`/�STMk/�/"D�/�-O/�/�H�/�?�'?�/�/i?�GIFs?�?�%�?F?X?�?�JPG�?!O�%`O�?�?qO�
JS{OĤO��7C�OOO%
�JavaScri3pt�O�?CS�O(_��&_�O %Ca�scading �Style Sh�eetsT_��
A�RGNAME.D)T�_��� \�_U_зA�T�_�_�PDI'SP*�_���To��_�QNa\oo
TP�EINS.XML��o�_:\�o]o�QC�ustom To�olbar�oiPASSWORDSo~��FRS:\#��oD`Passwo�rd Configd���<�� ��+�=��a���� ��&���J�ߏn���� ��9�ȏ2�o�����"� ��ɟX��|��#��� G�֟k������0�ů T����������C�U� �y������>�ӿb� ������-ϼ�Q��J� ��ϫ�:�����p�� ��)�;���_��σ�� $߹�H���l����� 7���[�m��ߑ� �� ��V���z�����E� ��i���b���.���R� ��������AS�� w�*<�`� ��+�O�s� �8��n/� '/��]/��//z/ �/F/�/j/�/?�/5? �/Y?k?�/�??�?B? T?�?x?O�?OCO�? gO�?�O�O,O�OPO�O �O�O_�O?_�O�Ou_ _�_(_�_�_^_�_�_ o)o�_Mo�_qo�oo �o6o�oZolo�o% �o[�o�� D�h���3�� W��������@��� �v����/�A�Џe� 􏉟��*���N��r��������$FIL�E_DGBCK �1V������ < ��)
SUMMA�RY.DG#�Ϝ�MD:W���ې�Diag Sum�mary����
C?ONSLOG��p����ۯ���Con�sole log����	TPACC�N�v�%^������TP Accou�ntin=���F�R6:IPKDM�P.ZIPϿӘ
�� ϧ���Exception$�ջ���MEMCHECKБ�������/�Me�mory Dat�a����l�)��RIPE��ϒ��'߶�%�� Packet L<����L�$�e���S�TAT!��߯�� %C�Sta�tus��`�	FTAP������1��mment TB�D4�`� >I)ETHERNEy���f�w�瑱Et�hernL�3�fi�guraCϫ��DCSVRF(�� ��9����� verify all<����M.c��DIFF1��)���=�S�diff��t�f���CHG01������`C����kv�- 	29 2���hz�3���K ��rVTR�NDIAG.LS�w(:���� �Ope��N� ��n�ostic����)VDEV�DAT�������Vis�Dev�ice�+IMG@��./@/�/<�k$�Imagw/+U�P ES/�/FORS:\?\=���Updates OList\?��� �FLEXEVEN���/�/�?���1 ?UIF EvO�O����,�t)
P�SRBWLD.C	MOϜG2#O^?0��PS_ROBOW�ELU���:GIG��ϾO�?�O��Gi�gE�(O��N�A��)�AHADO�W�O�O�Oi_��S�hadow Ch�ange����a��)RRCMERR�a_F_X_�_���PC�FG Error�q tail�_ M�A�m�CMSGLIB�_�_�_so�B�6e��|0ico+a7�)_`ZD�O�o�\o�o��ZDPa�d�o l )RNO�TI��o�ow��Notific�� F�AG���՟ ����(���L��p� �����5�ʏ܏k� � ��$�6�ŏZ��~�� ����C�؟g������ 2���V�h�������� ¯Q��u�
����@� ϯd�󯈿��)���M� �����ϧ�<�N�ݿ r�ϖ�%ϣ���[��� ��&ߵ�J���n߀� ߤ�3�����i��ߍ� "��/�X���|��� ��A���e������0� ��T�f�������=� ����s���,>�� b����'�K� ���:�Gp ��#��Y�} /$/�H/�l/~// �/1/�/U/�/�/�/ ? �/D?V?�/z?	?�?�? ??�?c?�?
O�?.O�? RO�?_O�OO�O;O�O �OqO_�O*_<_�O`_ �O�_�_%_�_I_�_m_ �_o�_8o�_\ono�_ �o!o�o�oWo�o{o "�oF�oj�ow� /�S����� B�T��x������=��ҏa������,����$FILE_FR�SPRT  ��������A�MDONL�Y 1VU��� 
 �)MD�:_VDAEXTP.ZZZ3�䏻��ʛ6%NO� Back fi�le ���S�6)�����@�	�M�v� ����)���Я_����� �*���N�ݯr���� ��7�̿[�ٿϑ�&� ��J�\�뿀�Ϥ϶� E���i���ߟ�4��� X���eߎ�߲�A��� ��w���0�B���f���ߊ��E�VISB�CKs�]���*.�VD����U�FR�:\��ION\DOATA\��w�U��Vision VD��!�[�m��� ��{��D�����z� ��3E��i��� .�R���� A�Rw�*� �`��/��O/ �s/�/@/�/8/�/\/ �/?�/'?�/K?]?�/��??�?4?F?�?;�L�UI_CONFIoG WU���>�; $ �3x�{U�=OOOaOsO�O�O�I%@|x�?�O�O�O __'\�OJ_\_n_�_ �_)_�_�_�_�_�_o �_4oFoXojo|o�o%o �o�o�o�o�o�o0 BTfx�!�� �����,�>�P� b�t��������Ώ�� ����(�:�L�^�p� �������ʟܟ� ��$�6�H�Z�l���� ����Ưدꯁ�� � 2�D�V�h��������� ¿Կ�}�
��.�@� R�d����ϚϬϾ��� ��y���*�<�N�`� �τߖߨߺ�����u� ��&�8�J���[�� ������_������ "�4�F���j�|����� ����[�����0 B��fx���� W��,>� bt����S� �//(/:/�^/p/ �/�/�/=/�/�/�/ ? ?$?�/H?Z?l?~?�? �?9?�?�?�?�?O O �?DOVOhOzO�O�O5O �O�O�O�O
__�O@_ R_d_v_�_�_1_�_�_ �_�_oo�_<oNo`oPro�o�o&h�`x�o��c�$FLUI_�DATA X�����a�)a�dRESUL�T 2Y�ep� �T�/w�izard/gu�ided/ste�ps/Expert�o?Qcu�����������Skip Gpa�nce and �Finish Setup�D�V�h� z�������ԏ����&h �`.)`|�e!�0 �2`�!��c�aA��ps�������ԟ� ��
��.�@�R��2o y���������ӯ��� 	��-�?�Q�)e�)c�A�3�E�W�g�rip*pu�ۿ����#� 5�G�Y�k�}Ϗϡ�`� ����������1�C� U�g�yߋߝ�\�n�����ߤ�b�g�%pTi�meUS/DST ��?�Q�c�u������������
�Enable��(�:�L� ^�p��������������� �b�a����0�����#�24*� ������ 1C��y��� ����	//-/?/ Q/"4F\�$q?RegionT/�/ �/??+?=?O?a?s?��?�?�AmericaϿ�?�?�?O O+O=OOOaOsO�O�O�)aym//�O�/�/>#sditor�O7_ I_[_m__�_�_�_�_��_�_� Touc�h Panel � S (recommenp)�_>oPo boto�o�o�o�o�o�o�o�L��O�O5�O	_>Racces�?� ���������,�>���Conn�ect to N?etworkM��� ������̏ޏ����P&�8�J��H�^ 9�+=S!_PIntroduct�/ �����*�<�N�`� r������Ϻ�̯ޯ� ��&�8�J�\�n������� ��w�����|YVSafet�A $�6�H�Z�l�~ϐϢ� �������ϩ�� �2� D�V�h�zߌߞ߰��� �����߷�ɿ��[ �k�}�������� ������1�C��g� y��������������� 	-?[(�5��-�Q��� ��"4FXj |�M������ //0/B/T/f/x/�/ �/[m�/�?? ,?>?P?b?t?�?�?�? �?�?�?��?O(O:O LO^OpO�O�O�O�O�O �O�O�/_�/3_�/Z_ l_~_�_�_�_�_�_�_ �_o o2oDoU_hozo �o�o�o�o�o�o�o
 .@�Oa#_�G_ �������*� <�N�`�r�����Uo�� ̏ޏ����&�8�J� \�n�����Q��uן ����"�4�F�X�j� |�������į֯诧� ��0�B�T�f�x��� ������ҿ俣��ǟ )�;���b�tφϘϪ� ����������(�:� ��^�p߂ߔߦ߸��� ���� ��$�6���?� �c��Oϴ������� ��� �2�D�V�h�z� ��K߰���������
 .@Rdv�G� ��k����* <N`r���� ����//&/8/J/ \/n/�/�/�/�/�/�/ ����1?�X?j? |?�?�?�?�?�?�?�? OO0O�TOfOxO�O �O�O�O�O�O�O__ ,_>_�/?!?�_E?�_ �_�_�_�_oo(o:o Lo^opo�oAO�o�o�o �o�o $6HZ l~�O_a_s_��_ �� �2�D�V�h�z� ������ԏ�o�
� �.�@�R�d�v����� ����П⟡��'� �N�`�r��������� ̯ޯ���&�8�I� \�n���������ȿڿ ����"�4��U�� y�;��ϲ��������� ��0�B�T�f�xߊ� I������������� ,�>�P�b�t��Eϧ� i���Ϗ���(�:� L�^�p����������� ���� $6HZ l~������� ���/��Vhz �������
/ /./��R/d/v/�/�/ �/�/�/�/�/??*? �3W?�?C�?�? �?�?�?OO&O8OJO \OnO�O?/�O�O�O�O �O�O_"_4_F_X_j_ |_;?�?_?�_�_�?�_ oo0oBoTofoxo�o �o�o�o�o�O�o ,>Pbt��� ���_�_�_�_%��_ L�^�p���������ʏ ܏� ��$��oH�Z� l�~�������Ɵ؟� ��� �2����w� 9�����¯ԯ���
� �.�@�R�d�v�5��� ����п�����*� <�N�`�rτ�C�U�g� �ϋ�����&�8�J� \�n߀ߒߤ߶��߇� �����"�4�F�X�j� |����������� �����B�T�f�x��� ������������ ,=�Pbt��� ����(�� I�m/����� �� //$/6/H/Z/ l/~/=�/�/�/�/�/ �/? ?2?D?V?h?z? 9�?]�?��?�?
O O.O@OROdOvO�O�O �O�O�O�/�O__*_ <_N_`_r_�_�_�_�_ �_�?�_�?o#o�OJo \ono�o�o�o�o�o�o �o�o"�OFXj |������� ���_'ooK�u�7o ������ҏ����� ,�>�P�b�t�3���� ��Ο�����(�:� L�^�p�/�y�S���ǯ ��� ��$�6�H�Z� l�~�������ƿ��� ��� �2�D�V�h�z� �Ϟϰ��ρ������� �ۯ@�R�d�v߈ߚ� �߾���������׿ <�N�`�r����� ��������&����� 	�k�-ߒ��������� ����"4FXj )������� 0BTfx7� I�[�����// ,/>/P/b/t/�/�/�/ �/{�/�/??(?:? L?^?p?�?�?�?�?�? ��?�O�6OHOZO lO~O�O�O�O�O�O�O �O_ _1OD_V_h_z_ �_�_�_�_�_�_�_
o o�?=o�?ao#O�o�o �o�o�o�o�o* <N`r1_��� �����&�8�J� \�n�-o��Qo��uow� ����"�4�F�X�j� |�������ğ���� ��0�B�T�f�x��� �������ᯣ��� ۟>�P�b�t������� ��ο����՟:� L�^�pςϔϦϸ��� ���� ��ѯ���?� i�+��ߢߴ������� ��� �2�D�V�h�'� ������������
� �.�@�R�d�#�m�G� ����}�����* <N`r���� y���&8J \n����u��� ����/��4/F/X/j/ |/�/�/�/�/�/�/�/ ?�0?B?T?f?x?�? �?�?�?�?�?�?OO ���_O!/�O�O�O �O�O�O�O__(_:_ L_^_?�_�_�_�_�_ �_�_ oo$o6oHoZo lo+O=OOO�osO�o�o �o 2DVhz ���o_���
� �.�@�R�d�v����� ����}oߏ�o��o*� <�N�`�r��������� ̟ޟ���%�8�J� \�n���������ȯگ ����Ϗ1��U�� |�������Ŀֿ��� ��0�B�T�f�%��� �Ϯ����������� ,�>�P�b�!���E��� i�k�������(�:� L�^�p�����w� ���� ��$�6�H�Z� l�~�������s����� ����2DVhz �������
 ��.@Rdv�� �����/�� ��3/]/�/�/�/�/ �/�/�/??&?8?J? \?�?�?�?�?�?�? �?�?O"O4OFOXO/ a/;/�O�Oq/�O�O�O __0_B_T_f_x_�_ �_�_m?�_�_�_oo ,o>oPoboto�o�o�o iO{O�O�O�O(: L^p����� �� ��_$�6�H�Z� l�~�������Ə؏� ����o�o�oS�z� ������ԟ���
� �.�@�R��v����� ����Я�����*� <�N�`��1�C���g� ̿޿���&�8�J� \�nπϒϤ�c����� �����"�4�F�X�j� |ߎߠ߲�q��ߕ��� ���0�B�T�f�x�� ������������� ,�>�P�b�t������� ����������%�� I�p����� �� $6HZ �~������ �/ /2/D/V/w/ 9�/]_/�/�/�/
? ?.?@?R?d?v?�?�? �?k�?�?�?OO*O <ONO`OrO�O�O�Og/ �O�/�O�O�?&_8_J_ \_n_�_�_�_�_�_�_ �_�_�?"o4oFoXojo |o�o�o�o�o�o�o�o �O_�O'Q_x� �������� ,�>�P�ot������� ��Ώ�����(�:� L�U/y���eʟ ܟ� ��$�6�H�Z� l�~�����a�Ưد� ��� �2�D�V�h�z� ����]�o��������� �.�@�R�d�vψϚ� �Ͼ������ϳ��*� <�N�`�r߄ߖߨߺ� ���������ӿ�G� 	�n��������� �����"�4�F��j� |��������������� 0BT�%�7� �[����� ,>Pbt��W� ����//(/:/ L/^/p/�/�/�/e�/ ��/�?$?6?H?Z? l?~?�?�?�?�?�?�? �?? O2ODOVOhOzO �O�O�O�O�O�O�O�/ _�/=_�/d_v_�_�_ �_�_�_�_�_oo*o <oNoOro�o�o�o�o �o�o�o&8J 	_k-_�Q_S�� ���"�4�F�X�j� |�����_oď֏��� ��0�B�T�f�x��� ��[���󟷏� ,�>�P�b�t������� ��ί�򯱏�(�:� L�^�p���������ʿ ܿ���џ�E�� l�~ϐϢϴ������� ��� �2�D��h�z� �ߞ߰���������
� �.�@���I�#�m�� YϾ���������*� <�N�`�r�����Uߺ� ������&8J \n��Q�c�u�� ���"4FXj |�������� //0/B/T/f/x/�/ �/�/�/�/�/�/�� �;?�b?t?�?�?�? �?�?�?�?OO(O:O �^OpO�O�O�O�O�O �O�O __$_6_H_? ?+?�_O?�_�_�_�_ �_o o2oDoVohozo �oKO�o�o�o�o�o
 .@Rdv�� Y_�}_��_��*� <�N�`�r��������� ̏ޏ����&�8�J� \�n���������ȟڟ 쟫��1��X�j� |�������į֯��� ��0�B��f�x��� ������ҿ����� ,�>���_�!���E�G� ����������(�:� L�^�p߂ߔ�S����� ���� ��$�6�H�Z� l�~��Oϱ�s����� ��� �2�D�V�h�z� ��������������
 .@Rdv�� ���������� 9��`r���� ���//&/8/�� \/n/�/�/�/�/�/�/ �/�/?"?4?�= a?�?M�?�?�?�?�? OO0OBOTOfOxO�O I/�O�O�O�O�O__ ,_>_P_b_t_�_E?W? i?{?�_�?oo(o:o Lo^opo�o�o�o�o�o �o�O $6HZ l~������ �_�_�_/��_V�h�z� ������ԏ���
� �.��oR�d�v����� ����П�����*� <������C����� ̯ޯ���&�8�J� \�n���?�����ȿڿ ����"�4�F�X�j� |ώ�M���q��ϕ��� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t���� ����������%��� L�^�p����������� ���� $6��Z l~������ � 2��S�w 9�;�����
/ /./@/R/d/v/�/G �/�/�/�/�/??*? <?N?`?r?�?C�?g �?�?�/OO&O8OJO \OnO�O�O�O�O�O�O �/�O_"_4_F_X_j_ |_�_�_�_�_�_�?�? �?o-o�?Tofoxo�o �o�o�o�o�o�o ,�OPbt��� ������(��_ 1ooU��Ao����ʏ ܏� ��$�6�H�Z� l�~�=����Ɵ؟� ��� �2�D�V�h�z� 9�K�]�o�ѯ����
� �.�@�R�d�v����� ����п������*� <�N�`�rτϖϨϺ� ���ϝ�����#��J� \�n߀ߒߤ߶����� �����"��F�X�j� |������������ ��0�����u�7� ������������ ,>Pbt3�� ����(: L^p�A��e�� ��� //$/6/H/Z/ l/~/�/�/�/�/�/� �/? ?2?D?V?h?z? �?�?�?�?�?��?� O�@OROdOvO�O�O �O�O�O�O�O__*_ �/N_`_r_�_�_�_�_ �_�_�_oo&o�?Go 	Oko-O/o�o�o�o�o �o�o"4FXj |;_������ ��0�B�T�f�x�7o ��[o��Ϗ����� ,�>�P�b�t������� ��Ο����(�:� L�^�p���������ʯ ��ӏ����!��H�Z� l�~�������ƿؿ� ��� �ߟD�V�h�z� �Ϟϰ���������
� �ۯ%���I�s�5��� �߾���������*� <�N�`�r�1ϖ��� ��������&�8�J� \�n�-�?�Q�c����� ����"4FXj |�������� 0BTfx� ����������/ ��>/P/b/t/�/�/�/ �/�/�/�/??�:? L?^?p?�?�?�?�?�? �?�? OO$O��/ iO+/�O�O�O�O�O�O �O_ _2_D_V_h_'? y_�_�_�_�_�_�_
o o.o@oRodovo5O�o YO�o}O�o�o* <N`r���� ��o���&�8�J� \�n���������ȏ�o 鏫o��o4�F�X�j� |�������ğ֟��� ���B�T�f�x��� ������ү����� ُ;���_�!�#����� ��ο����(�:� L�^�p�/��Ϧϸ��� ���� ��$�6�H�Z� l�+���O����߇��� ��� �2�D�V�h�z� �����������
� �.�@�R�d�v����� ����}��ߡ����� <N`r���� �����8J \n������ ��/����=/g/ )�/�/�/�/�/�/�/ ??0?B?T?f?%�? �?�?�?�?�?�?OO ,O>OPObO!/3/E/W/ �O{/�O�O__(_:_ L_^_p_�_�_�_�_w? �_�_ oo$o6oHoZo lo~o�o�o�o�o�O�O �O�O2DVhz �������
� �_.�@�R�d�v����� ����Џ�����o �o�o]��������� ̟ޟ���&�8�J� \��m�������ȯگ ����"�4�F�X�j� )���M���q�ֿ��� ��0�B�T�f�xϊ� �Ϯ���ѿ������ ,�>�P�b�t߆ߘߪ� ��{��ߟ��ÿ(�:� L�^�p������� ���� ����6�H�Z� l�~������������� ����/��S� �������
 .@Rd#��� �����//*/ </N/`/�/C�/�/ {�/�/??&?8?J? \?n?�?�?�?�?u�? �?�?O"O4OFOXOjO |O�O�O�Oq/�/�/�O 	_�/0_B_T_f_x_�_ �_�_�_�_�_�_o�? ,o>oPoboto�o�o�o �o�o�o�o�O_�O 1[_����� �� ��$�6�H�Z� o~�������Ə؏� ��� �2�D�V�' 9K��oԟ���
� �.�@�R�d�v����� ��k�Я�����*� <�N�`�r��������� y���������&�8�J� \�nπϒϤ϶����� ���Ͻ�"�4�F�X�j� |ߎߠ߲��������� �˿ݿ�Q��x�� ������������� ,�>�P��a������� ��������(: L^�A�e�� �� $6HZ l~������ �/ /2/D/V/h/z/ �/�/�/o�/��/� ?.?@?R?d?v?�?�? �?�?�?�?�?O�*O <ONO`OrO�O�O�O�O �O�O�O_�/#_�/G_ 	?_�_�_�_�_�_�_ �_�_o"o4oFoXoO |o�o�o�o�o�o�o�o 0BT_u7_ ��oo����� ,�>�P�b�t������� ioΏ�����(�:� L�^�p�������e� �ӟ���$�6�H�Z� l�~�������Ưد� ���� �2�D�V�h�z� ������¿Կ����� �۟%�O��vψϚ� �Ͼ���������*� <�N��r߄ߖߨߺ� ��������&�8�J� 	��-�?ϡ�c����� �����"�4�F�X�j� |�����_��������� 0BTfx����m�������$FMR2_GR�P 1Z��� �C4�  B��	 ��;M8E��� F@ c�5�Wo�
8J��N�Jk�I'PK�Hu��IP�s�F!��{?� � ��89�<�9�89�6C'6<,�5��{A� � /+BH5B�x10 !@�33;"�33�7]/n-^8@UUT�*@9 �� {��>u.�>*��<���{�>���>��l�=<��=�U��=�v!>1
�{:�ܜ:2B�8'Ŭ9I�R7���9f�͛/$?o/!?Z?E?~?�i?�?��_CFG� [T �?�? OO�;NO {
F0HA� M@�<RM_CHKTYP  ��&(� ROM�c@_MINi@������@�T XS�SB�3\� 9�O���C��O�O�5TP_DEWF_Oz��&>	WIRCOMh@_��$GENOVR/D_DO�F��G]�THR�F ddUd�MT_ENB9_ ^MPRAVC]�G��@ �[F�@ G��@GA�w\H͊#Iv0�Iά �?�O�o�o(oK* ��QOUc�PAKRK< �@��oIo�o�o�o��?C�  D�o�ht1A|A$ B�L�.rN�i�O�PSMT�d�Y*�@t�$�HOSTC�21e��@���7 kMC��T{����  27.0z2�1�  e� _�q�������M�Ə؏���������	anonymous#� Q�c�u��������6�������F�'� 9�K�]�o��������� ɯ쟆�0��#�5�G� Y�k�����ҟ���׿ �����1����g� yϋϝ���������� 	��-�p��ϔ����� ��ܿ���������H� )�;�M�_�q������ ���������D�V�h� z�|�R��ߑ������� �����!3Eh� �������� *�<�N�PA��ew ��������/ /<n3/a/s/�/�/ �/���/$/?X 9?K?]?o?�?��?�? �?�?�/�?B/#O5OGO YOkO}O�/�/�/�O�? �O,?__1_C_�?g_ y_�_�_�_�OT_O�_�	oo-o?o�~�qEN�T 1f�y� � P!�_�o  �p~o�o�o�o�o �o'�o3\�D �h������ �G�
�k�.���R��� v���鏬��Џ1�� U��N���z���r�ӟ �������ޟ,�Q�� u�8���\�����ᯤ�����گ;���_�"�?QUICC0l�H�Z���~�1��������~�2����[�!?ROUTER\�8��Jϫ�!PCJO�G�χ�!19�2.168.0.�10��z�CAMP�RT����!��1��#�
�RTu�'�9���� !Soft�ware Ope�rator Pa�nelw�����`dN�AME !mj!�ROBO���S_CFG 1emi� �A�uto-star�ted�DFTP�O���O�_���O�� ������c_>�P�b� t����+��������� �@\�n��a�� ��x������ '9Kn��� �����O�O�O�O V,/�k/}/�/�/�/ v�/�/�/??B/�/ U?g?y?�?�?�?�/ /(/*?O^/?OQOcO uO�OJ?�O�O�O�O�O O�O)_;_M___q_�_ �?�?�?�_�O�_2Oo %o7oIo[o_o�o�o �o�_�olo�o!3 EW�_�_�_��o� o�����oA�S� e�w����.���я� ����\n��s� �������͟ߟ񟴏 �'�9�K�]������ ����ɯۯ�0�B�T� f�h�Y���}������� ſ�������1�T� ֿg�yϋϝϯ�����_ERR g������PDUSIZW  V�^t�����>	�WRD ?�J�7��  guestVƀI�[�m�ߑߣ���S�CDMNGRP �2hJ���C�7�V�8V�K��� 	P01.0�3 8�   �e�?��  �;  �  �� ���ߛ����@�-��������x����0���y�d������,�>�P���~��  D��d����������_�GROU��i��J����	���5{��QUP�3��������TYC �����TTP_AUT�H 1j�� <�!iPenda�n��%`Ϗ�!�KAREL:*8%.@KCUe�wM VISION SET����V�K��J( @:�^p������CTRL �k����%V�
D�K�FFF9E3��5�FRS:D�EFAULT3,�FANUC W�eb Server3*! 5���1�C����/�/�/�/�/?��W�R_CONFIGw l�� 3/���IDL_CPU�_PCR V�B��8�u0 BH[5MI�Nf<!�y5GNR_�IO���V���]0N�PT_SIM_D�O�6�;STAL�_SCRN�6 ����INTPMOD�NTOL�7�;�!R�TY�8u1�6� ��E�NB�7��Y4OL_NK 1m��E� }O�O�O�O�O�O�OaBMASTE�0��aB�SLAVE n���URAMCAC�HE_�2O��O_�CFGI_`CaSUO���l_]RCMT_O�PR �2�ʟSYCL�H_{UL _ASG s1o��#�
 �O o o2oDoVohozo�o �o�o�o�o�o�o�K�RWNUM���
]R�IPF_XWRTRY_CN�_{U�1��ӊ|A��� ]R�PfR�p'^=з=�]0P_�MEMBERS �2q��� $�%�r����w��]0�RCA_ACC �2r��  V��# 
�� �/� 3y  5Ө�(�� S�5`��H�c�U�  �V�5�BUF00�1 2s��= ��u0  u0[�փބބ�#ބ-?�  ?��	�փ

���+�;�L�[��m�|�������������Z��փ~�~�U!~�1~�B~�Q~��c~�r~��u0(� M�u0��`x�u0I_�+��~��~���u0�s8}րuփ�,��Cu0$�QYu04�o@�%��4փ�E&�T&�=�6�w>pE� r0��ք ք/�ք����bքq�ք�ք�ք�ք�Jք�ք�փ��2�� ҃ց܁ց�������k(
�� ���ց���� ��%��-��5�� =��E��M��U�� ]��e��m��u�� }�ց������������ ���������������� ����Ő��͐��Ր�� ݐ��吉��ց���� �����������ցx���$�_@�,��!�5�!�F�D�t(L�N�T��]��e� ᢮�t��}�ᢅ����q�`��ᢝ� ᢥ�᢭�ᢵ�ց��3ɯ҅�^"��^" ��` ��8���"� #�"%�3�"5�C�" E�S�"U�c�"e�s� "u���&񄓓��ҕ� ���ҥ����ҵ�ó�� Ő��͐��Ր��ݒ� ���&�������� ���&��+�*�-� ;�*�O�D��M�[��� ]�k��·�t����� �������¥�����X����gQ2t��4,%&�&�<&�K���25�HIS��v�� �S� 2�023-07-2���Y"{O�q8 U�p����������������V�Y&E�19Q�|B;��p:m�L^p���p����s!8Q�,>Pbtd�Y!�Y!׀���ҫ�s!�:�s
��7��q� /"/4/F/X/j/|/�/ �/���/�/�/?? 0?B?T?f?x?�/�/�? �?�?�?�?OO,O>O PO�?�?�O�O�O�O�O �O�O__(_z#�ȠP/�A�e�:- dU��Qc3_�_�_�_�_�_�oo1>  dA �d0oo�o�o�o �o�o�o�o��|_E�Wi{���� �c�io��r�- ' L�z�^iO{O �/�A�S�e�w����� ����eO�����+� =�O�a�s�����Ώ�� ��ߟ���'�9�K� ]�o�����ʟ��ɯۯ ����#�5�G�5_"� ��T_f_0e�ӹ� ƿؿ���� �2�D�h2oDoVh"� U� �ϲ����������� 0���f�xߊߜ߮� ���ߛ- ��߼-  �- �����B�T� f�x���������� �-��,�>�P�b�t� ������������� (:L^p�� �������� $�6HZlZ�l�I_�CFG 2wz�� H
Cycl�e Time��Busy�Idyl��min}=�Up���Read�gDow�� �}�Count��	Num ���ȩ`,S�7!EQPR�OG�xz����p/�/�/�/�/�/�?�@USDT_ISOLC  z����pJ23_�DSP_ENB � B;�c0INC� ys=S�P0A �  ?�  =�?��<#�
O1�9:�o �1�?�?�S��?O\7OB� C�l3��6"AG_GROUP 1zB;;�r<� �3(�	nOO?��/�OS�Q�O�O�O_�O0_�B_T_f_��?IG�_IN_AUTO�/D�:c0POSRE�*O<FKANJI_�MASK�V�ZKA�RELMON {z�h/S�y+_DoVo@hozo�o�b�#|�'�~3S��e�_4K�CL_L�PNUM�p0�o$KEYLO�GGING�`����q{5� LANGU�AGE z��Jp�DEFA�ULT Xqh�LGf�}�*��Sѽx�0�  R��H  �S�'�� + �SЛS�?)7�;��
�q(U�T1:\�o�  ����0�=�O�a�x�������(3o�c��LN_DISP �~�?��O�O��O�CTOL9�S�Dz�� K1�1O�GBOO	Kq0i}d���������X�|����ϟៀ���us�'��	m��yjA%;o�?�1�k�_BUFF 2��B; �S�2 �����*2ү�� � -�$�6�c�Z�l����� ��Ͽƿؿ���)� ��2�_π3��DCS ��)�2�1$�c������������v�IOw 2��� �3�jA�6�F�X�j� ~ߎߠ߲��������� ��0�B�V�f�x�������������ER/_ITM?>d�_?� Q�c�u����������� ����);M_�q���I��SE�V�`s=�TYP?>.�!3��Q�RSTt�SCRN_FL 2��� ��ϧ���0�//DTPp??��C�NGNAMpl4��Jrr�UPS�SGI\�U{5�!�_LOAD'@G �%@*%DMA�Yɥ�/G�MAXU�ALRM�b�QC���{5
�"�!_PRD�$�P a�%�� C��i�ٯè)3H@�P 2�w� �ZƦ	O!t�0��0�P?���2�?�?�?�? ���?+OOOO2ODO�O pO�O�O�O�O�O_�O '_
__]_H_�_l_�_ �_�_�_�_�_�_�_5o  oYoDo}o�oro�o�o �o�o�o�o1U gJ�v���� �	��-�?�"�c�N� ��j�|������̏� ���;�&�_�B�T��� ������ݟ�ҟ����7��'DBGDEF �25?1>1@�R��_LDXDISA�m ?+�MEMO_{APg E ?@+
 d����ү������,�>�� F�RQ_CFG ��27h�A �@i���!�<?4d%A�Э�R�d�z2�2;��4*��/�� **:�!��� ȟ�!�,�>�k�b�t� �ϘϪ���#�25 ���`��'�� �6�,(�� ~���lߩߐ��ߴ��� ���'��K�]�D���h�������*IS�C 1�@)� � )�#��4i�9�$�r�]��������_MSTR� ����SCD 1�������� ,P;t_q� �����& L7p[��� ���/�6/!/Z/ E/~/i/�/�/�/�/�/ �/�/ ??D?/?A?z? e?�?�?�?�?�?�?�? OO@O+OdOOO�OsO �O�O�O�O�O_�O*_ _N_9_^_�_o_�_�_��_�_�_�_o��MK�g������&o$M�LTARMf��:۷Qb �b���o�dQ�METPU܋�b����ND�SP_ADCOLx�ef��nCMNT�o �eFN�`�o�gFSTLIw�� ���g~�c��|�t�ePOSCF5w=�nPRPM�o�y�ST�`1��� 4��#�
��� �!��!�#�5�w�Y� k��������ŏ׏� ���O�1�C���o��a�SING_CHK�  $MODAe���OkQn���DEV 	��	�MC:�HSI�ZE��`ȿ�TA�SK %��%$�12345678�9 `�r���TRI�G 1��� l Q�����Lٮ��L�B��YP-�L�Ք��E�M_INF 1��ۻ`)AT?&FV0E0��k��)S�E0V1&�A3&B1&D2�&S0&C1S0}=Z�)ATZk�����Hÿ�z�߯���A�C���g�Nϋ��� Q���u������� �Ͽ@�w�d�v�)Ϛ� U߾��߷��ߧϹ�*� �����r�}�7ߨ��� �������&��J� \���3�E�W�i��� ����5�4��X |�u�e�w���� ����0B��f�� EO�{��// �>/�'�/K �/�//�/�?�/'?�L?3?p?�NITO�RPpG ?�  � 	EXEC�1c�22�83�84��85�8���67�88
�89c�2:"D�2 D�2D�2D�2D�2 D�2D BDBDB�C2%H21H2=H2�IH2UH2aH2mH2�yH2�H2�H3%H3�1H3�2��R_GRP_SV 1�@�� (w���<�� ��>%���6����u�=���J�_D�20�ySION_D�Bɐ�͝a  ��`�☾T �Z`��W��ps�>f0N   #v�W�G�-ud1��/oAoSo�aPL_NAME !Q��|`�!Def�ault Per�sonality� (from FsD)�P�bRR27Q� 1�L�XL��x|a�P dzr�o�o�o�o# 5GYk}��� ������1�C���2�on���������@ȏڏ������<]� :�L�^�p���������@ʟܟ� �[i*�)�":�
)�^�]dPM��� ������ү����� ,�>�P�b�t�����g� y�ο����(�:� L�^�pςϔϦϸ��� �ϫ����$�6�H�Z� l�~ߐߢߴ����������� �2� F�@ G&h G�]gSP  �_�q�]bd[�C���� ������D�7�Zj��	�p��=�@� -� X�N�`�r����������SP�0��	]b-�	�`B�<N`:�oA�b����? A�  �	W�kV]`�S ]`���PCT���P�h�`)  �  u$�T&"� C�gyd���:\kR6R 1�ti�P�*0 � �f2|`  @D��  !?�#X�,?]`!]aA/���%iJ-;�	�l,"	 �߀pJn ��NP`e  � � w� �� � ��"�SPK�K ���K=*�J����J���J9�٧�U�p��/SP@�_f��"j�@��(E14!�/�#�N����;f,1��� �a�������-�@¾ - T1�HZ0Z0� ��/  >c�=���>�Q ���o���l? �?��2-!�3�&. Up�Pm P� ��P_�  ��P�F��*O�%	'� �� HBI� ��  ���&:��ÈlOÈ=�s�̈́E�"@�O@�@�>!�O/K"���&&�&�Q_  '�`.T�!-0@2��O@����"=0@A?�C� C�PC��� Ca0Ce0Ci=�%��A�% 0� �Pl�-_hhX�'B�P��Q���A�U]aDz �on?3ooCoio�O��dIA�R�TZ��A����  �4@?��ff���o�ono  #{�!8�@9GzC>L�@�0(!�*(�@ uu�0�v�i{!t#t$�C�?]t�@,��<
6�b<߈;܍��<�ê<���<�^¬/�C�A�K"�#,"� �?fff?�@?&�&���@�.8���J<?�\�D�N\��I�R!�-$�)% |�'��
�`$�oЏ�� �ߏ��<�'�`�r�0]����He�F| �� ҟ����m�����J���F�  F��~�BG�d GC�q V���R���ů���ԯ ���1��U�@��O�� �F�IG/�ӿ1���m� �0�B�T�:��o�{�33ϩ���ϸ������{An� ��_��EC��U��ϲ�d�?�؃ߊ��߮��Im�i4����C �CfPa0�¸�Ԑ0ؼ��@�@I���B�>�)A�C�A�IA��@?�?\����ú@ �������=q��A��Ay�I33@�0��@��C��1������(���C�����b��=q�Ů�����H��� G�� G��B�I��(E�ψ C�e�� I"�L�J�H�V@G5� E��x C��I3��J0�G��߀I�� 0 C ='�߀�k��������� ������"F1j Ug������ �0B-fQ� u�����/� ,//P/;/t/_/�/�/ �/�/�/�/�/??:? %?7?p?[?�??�?�? �?�? OO�?6O!OZO EO~OiO�O�O�O�O�O �O�O __D_/_h_z_�e_�_�_�_�_�_y�(΄�����r��<$e�U��o&o9�3�8�@oRo9я4Mgulo~o9Ѵ�VwQ�o�o4p�+4�]�m�i@�o(L:|u�P�r	P~~������_�0����{R��`G�2�W�}�h�  �`��ˏ���ڏ�����F�4�j�X� p�z��������ԟz����4�"�X�F�|����  2 F�@9�G&h�����9�B�&��)��C	�&�9�@-��9�o`�+�=�O��� ��{�Ħ�GAw\]�0����ɿ7�?��|p*9�t�9�9��9�{�
 ֿ9� K�]�oρϓϥϷ��π�������#�z�����hk�y��$�MR_CABLE� 2�hx i�ћqT�p@��¦�?>𦡆т����кƠ��C��ޱO8�tB�����8��ް.ޱF\�!�޶�ߕ��>���š��C�N�|�z����a}`r����	P��e����L�  ���C֠:��������a���!ްޱE�S "�4��ՠ�y�qBy�ԡ��HE����ls�޵;�aZ v�/ߘ���k������ C��L�>�8�f�\�n� ������������?��H�� oq<����ܸ���ܸ�*,** \�O�M �i������ Ël%% �2345678901i{ f��Rް�ް�ްޱ�
�not? sent 5��WpuTES�TFECSALG&#�egۺ�d.$���
>$���p�޴�޷Y/k/}/�/ �9UD1:\m�aintenances.xml�/��/  ��DEFAULTa�~\�GRP 2�M�  pė�޵ � �%1st �mechanic�al check,�ޱ�z3鰄1�?��[ph��?�?�?��?�?޲R3cont?rollerb4,O{?PO���?|O�O�O�O�OAMY=�O޲"8SްQ_��kG8_J_\_n_�_�JACO�__�_�6/_@oo(o:oLoBC[0�geW2. batteryPo�_�o��	�_�o�o�o�o_i�@dui@able  D50Pq��`���o������Addgre�as;޷f��-ް�#���{P�b��t�����A
ddoi0�/��+�?�� &�8�J�\�Adj7޶����<ް������
�؟���� �B#|too�����>ǟ�������ү�AO?verhau�Ow��"� xް,�3�:5��`�r��������ް$Q�пSV��  O�$�6�H�Z�lϻ��� ߿�Ϲ������ � 2߁�VߥϷ��Ϟ߰� ������5ߝ��k�� ��d�v�������� ��1��U�*�<�N�`� r������������� &8��\���� ��������M "q�X�|�� ���7I/m B/T/f/x/�/��/� /�/3/??,?>?P? �/t?�/�/�/�?�?�? �?OOe?:O�?�?�? �O�O�O�O�OO�O _ OO�OsOH_Z_l_~_�_ �O�_�__�_9_o o 2oDoVo�_zo�_�_�o �_�o�o�o
ko@ �o�ov�o���� �1�Ug<��`� r��������̏�-� �Q�&�8�J�\�n��� ����ȟ����� "�4���X�����˟�� ��į֯���I��m� ���f�x���������5��	 T¿�� �*�4�F�X�j�|ώ� �ϲ����������� 0�B�T�f�xߊߜ߮� ����������,�>�P�b�t����� � �b�?�  @�  ���	������H�Z�l��;*��** @�>� 7����������,>��e�^��� A���u��� EWi�Ugy� ����/�/ -/?/�/u/�/�/� �/�/�/??�/;?�M?_?�/�/����$MR_HIST� 2�>��0� �
 \
�$ 23�45678901P�?�4�?���?9� )O;O�?$O��O�O�O ^OpO�O�O_�O�O_ I_[___6_�_�_l_ �_�_�_o�_3o�_Wo io o�oDo�o�ozo�o��o�oA�d�0S�KCFMAP  ]>��08�ʡ1�`IYuON�REL  �5�rq�0[rEXCFENB�w
psXu�q�FNC��tJOG_OVLIM�wd�3\�[rKEY�w�=�_PAN�x+�\'�[rRUN �,��SFSPDTYPx�x�uZsSIGN�>�tT1MOT��q�[r_CE_GRoP 1�>�rs �2ڰ9���c��8��8 &�g����B�����x� 埜�ڟ�ҟ?�Q�� u�,�����b�ϯ��ȯ ���)�;�"�_�������|����7[qQZ_�EDIT��lw��T�COM_CFG 1�h}�u�&�8�� 
��_ARC_��r�5�yT_MN�_MODE�����yUAP_CPL�]��tNOCHEC�K ?h{ @ �������� ,�>�P�b�t߆ߘߪ������ߍ{NO_WAIT_L���ՀNT���h{w��c�2�_ERR߁2	�hy�1�6�����@*��q�����w�O`�}�g�| 
�����0��a<O�00 ?��5�O�5��p"�Y�PA�RAMa�h{��� ������1�� = O08 ZlHx���������.���R��ODRDSP�\ã��xOFFSET_CAR�bψ�DIS��S_A�w�ARK���OPEN_FILE��;��S�OPTION_IO!�3� �M_PRG %�hz%$*E/W.�WmO������00�%�d.2  �p�v� C�!	� ��h�!�f����hRG_DSBOL  �7rqK��?eRIENTT5O�p�aC��pqq�A fUT_SIM_D'or��h�VlLCT �@<�粛$;��9�ed`7�_PEX���4R[AT� d�u�4>�UP �q>�{ �OOOBOPI��$��2ރ�L��XL�x[3�0C�O�O�O�O �O�O__(_:_L_^_ p_�_�_�_�_�_�_�_ o�g2�O/oAoSoeo wo�o�o�o�o�oB�o �o1CUgy@�������f�o �~9@�!�N�P�K� ]�o���������ɏۏ ����#�5�G�Y�(� :�������şן��� ��1�C�U�g�y��� ��l�~�ӯ���	�� -�?�Q�c�u����������Ͽ�s�¯���  �2͠4A�!S�e�G� �ϓ���A��������������!�3� Q�W�uߗ���{ ��������	`����!�x�:�o@1?�Q��c�u�A�  ��V+��!+�21�� 9���s � h�p )  �  u$ �����)��&�_�J�Ѓ�^fBl@O�01����� �{D��0 ���$  �� @D� � ��?���X�,?+���+�D��������  ;��	l��	 ���pJ3 ������*  � �� � �I � ��Ou�H(��H3�k7HSM5G��22G���GN�3h��(ϙ�u�SCH50�R50������r�û�¾ 5 ��� �� �)���m�AK����+�²���801 io��p�u����� p �m3�P00� �  � ��u���q�	'� � �"I� � � ���o�=��q�1/C+�@Y/@_ Z�!�/��"������q�NA0�/  �'R0�$���CA0C���*C. ??\�q�p�Az
b0�lwhhXn�B� �1��~�p!�5��zn��?3�?�? O.OU/GD!N2K4a�+����@?�ff�ϏO�O3OC ���O�KA8+��OZ>LS ���J(+�:U�EV^I@9�9�#?"T� ,A<�
6b<߈;�܍�<�ê<���<�^�qd�_�AAp+���#|���?fff?p �?&�PD@�.��R�J<?�\�	bN\��U2�Q� @��Ao��`o�W%�O �o�o�o�o�o�o�o %7"[mD�|��,oNoPo���xF��  F��+�G�d GCFQ�T� �d���u�����ҏ�� ������/M��&
 ������2��������J��O�[�3 pޟw�b�������
B<�A3�墚?+�C������w�)�?�ؠH�O���s�
�4�-ț�C��C��ć�b��b�a��@I��	B>�)A��C�AIA���@�?�\������ú@ ����/��=q+�R!>��I33@0��@���C�1����[�����C���'��=�q�Ů���	H�� G��� G�B�I���(E�� C��^l��I"L�J��HV@G5�� E�x C����I3�J0��G���I��? E@� C�� E�0�i�Tߍߟߊ��� ���������/��,� e�P��t������ �����+��O�:�s� ^���������������  9$]oZ� ~������� 5 YD}h�� �����/
/C/ ./g/R/d/�/�/�/�/ �/�/	?�/-???*?c?�N?�?r?�?>�(I��3�^opR���5�5����?�?@�3ǭ8�OO@�4M�gu1OCO@��Vw�Q]OoO4p�+4�]�M�I�O�O�OP�O_�L:�P�RPC^>�_�l_�?x_�_�_�_�[R�_�_o�_XoBo-o  �@�Eo Wo�o{o�o�o�o_Q�0�o/{5?@uc���?��������A�O�  2 F@@ƷG&hl���@�Ba����ձC��@�@򯷏ɏۏ����"�@��oL�^�p�����@�?���AP@ŕ�d@�@�<���@�
 ����� "�4�F�X�j�|��������į֯�?ʶ����-K�y��$P�ARAM_MEN�U ?�E��  �DEFPULSE���	WAITT�MOUTL�RC�V_� SHE�LL_WRK.$�CUR_STYLvJ���OPT��N��PTB����C��R_DECSNW� 4U���%�N�I�[� mϖϑϣϵ����������&�!�SSREL?_ID  �E]Q��5�USE_PR_OG %0�%"���6�CCRc�G�]Q�8���_HOST !0�!���ߔ�ATTP���ӿ�����|4��_TIMEa��G֯�!�GDEB�UGE�0�6�GINP_FLMSK]���T�P���PGAʹ� |�;���CH����TYPE-�9�!��Q�z�u��� ����������
 )RM_q��� ����*%7 Irm������/��WORD �?	0�
 	�PRy��SMAI����RSUͱ=#T1E��S�	��J"�COL�Uf)�/��LVc� �@��`ȯ��dq�TRACEC�TL 1��E�:� AP% &�'AP;P�.�&D/T Q��E0� �D � �F;�+0̐10�[Q@92��92Ԑ92.3�56�Ȑ12f5/4/4	�/4
/4/4/2��=4�E4�M4�-4��54�e6/4/4�/4G�12/4/4./2� DDTp�	B��	B!D"D#�D$/13S���4��4�=4�E4��M4�-4�54�e4���4��4��4��4�S DEDD�D�12>3�E4� M4,?>?P?b?t?�?�? �?�?�?�?�?O�OC���	BWDS�T�PT�!XC�S�T�T�T��D�-f�E�E
FS�MT�UT0!XCVO hOzO�O�O�O�_�O�O �O
__._@_R_d_v_ �_�_�_�_�_�o�_o o*o<oNo`oro�o�o �o�o�o�o�&z '1KEo���������ɟ ۟����#�5�G�Y� k�}�������ůׯ� ����1�C�U�g�y� ��������ӿ���	� �-�?�Q�c�uχϙ� �Ͻ���������)� ;�M�_�q߃ߕߧ߹� ��������%�7�I� [�m��������� �����!�3�E�W�i� {�����k��������� %7I[m ������� !3EWi{�� �����//// A/S/e/w/�/�/�/�/ �/�/�/??+?=?O? a?s?�?�?�?�?�?�? �?OO'O9OKO]OoO �O�O�O�O�O�O�O�O _#_5_G_Y_k_}_�_ �_�_�_�_���_oo 1oCoUogoyo�o�o�o �o�o�o�o	-? Qcu����� ����)�;�M�_� q���������ˏݏ� ��%�7�I�[�m�� ������ǟٟ���� !�3�E�W�i�{����� ��ïկ�����/� A�S�e�w����������ѿ�����#��$�PGTRACEL�EN  "�  ��!���7�_UP �/���f�n�R��g�7�_CFG7 �f�P�!�g����ĭϸ�|I���  ����{�DEFSPD ���� �I���7�H_CONFI�G �f�N� U!�!�d-��F�  �0�P����LѶ!��7�IN~�T�RL ��ͦ�8l��a�PE����f���,Ѹ�7�WLIDù��	�ٿLLB 1��� �M�B<�B94�� M�%���Pպ� << �?�O�n�O� f���������� "���<�j�P�r�����8�������
Q��@3Ev��GRoP 1����"��@��
����!�AM�D�@ D�@ Cf� @ �1����	�	,�,����uG���F´F(BI pP:L�p�!��>�l7>�����/.� =�-=%�T/Q// N/�/r/�/�/0/�/�/�/?)??  DzN3W?!�
>??.?�? �?�?�?�?�?�?!OO EO0OBO{OfO�O�O�O��J)�A
V7.10beta1�� A��� R��!�A!��@?!{G�Q=y�#�B����$Q@�����B�l�4Q@�CA���QT �O�i_{_�_�_FTp�� �<��_�_�_�_.� � �O��O�0oBo,ofo�Po�o�A-�p��u0�mf��o��o����@�AWP�R�c Bf��B�>0uBHfs*�d!�!�PuMד��d����r�cx�tx����$|����0���<�-�@�F�0�A�3�3`�������KNOW_M  �"��ƾ��SV ��C�]�m? ��$��o�H�3�E�~�!����M���� �R	��ѐlb��^�~��hhXd��1q� (�0u8�4�,����MR�³��&��oj3������OADBANFWD�����ST�1 1�f��4�խY� !

��.�_�R�d�v� �������п�'�� �]�<�Nϓ�rτ����Ϻ����2����	��ݠ�<3���3 �/�A�S��4p߂��ߦ��5�������߂�6�(�:�L��7 i�{����8����X�����MA֠���b�OVLD � ��~�P�ARNUM  p�������SCHa� o�
����	�UPD����#b>b�_CMP_��d�����'�zER�_CHK���`�˒���RSu��ٯ��_MO֯�_��a�_RES_G
����
V_��ch �������/ 
/;/./_/R/d/7�DT�/9oУ/�/ �/;���/??;� !?@?E?;h�`??�? ;���?�?�?;��?x�?O;V 1��v|ߠ��@`}\�THR_INRu��f��dqFMASmS~O Z�GMN}O��CMON_QUEUE ����
��Qa�N U�N8�F�H SENDQ#�YEXE._UD B�E-P_ SOPTI�OW,PPROG�RAM %�J%�P<O��RTAS�K_Ic�u^OCFG ��O���_
`�DATA���k	P�
2ʕyo�o�o �o�olo�o�o	-��oQcu�:oIN+FO���Wm��DC ����(�:�L�^� p���������ʏ܏ ��$�6�H��w�t��Wl r)	a��K_�a�i�~��EN!Bd�ѹ�2Ԙ�Ga2̙� X�,		�=��=� ���@�N�9��$��8�8�`D��_EDIT �o�����dWERFL�OXdC�RGADJ7 �}�A���줁?
���AϦQ�������?�O  Bz��ga<8�
�v%$�\�èr-�fg�2���r	H�@mlocBBP����q@'�ǽ�*۰/ݲ **: �ֿ��q��.@A��ſ�K�@��c���\I)#Ⱥ��1�[ϩ�g�������w�A.@u�������O� ��K�5�/�A߻�e߷� �ߛ߭�'���#��� ��=��y�s���� ����������k��g� Q�K�]����������� ��C��?)#5� Y����� ��1�mg y������_/ 	/[/E/?/Q/�/u/�/ �/�/�/7?�/3??? )?�?M?�?�?�?�?{ȁ	&o0OŠOWOBD�t$ qO�KEO�OAO��O�O	�PREF S��ŠŠ
ϥ?IORITY�W��}�ӡMPDSP�Q��A�7WUT�V��Φ�ODUCT�Q�}��O��OGg�_�TG���R��vRHI?BIT_DO���[�TOENT 1��}� (!AF�_INEaPog�!tcpoGm�!ud6oon!�icm^o�vRX�Y��}��š)�� ��o�oŠ� �o�e�o:!^E W�{��������6�H�*uS����A�J�����£>�+��Ѷ�/��z���¤�r�}�A;�,  �P}�8��J�\�n�ť�߆Z@ߏ����ҟ�£]��ENHANCE S�i�}�A�dޏD�+�rV�D� _Sɡ�ӡPORT_N�UMbSŠ.U�ӡ_CARTRE��l	�SKSTyAaW�[SLGS`�ٸk�;�HPU�nothing L�)�;�M�]����������_�TEMP �څY���5q�_�a_seiban �OϯO(�N�9�r�]� �ρϺϥ�������� ��8�#�\�G߀�kߐ� �ߡ���������"�� F�1�C�|�g����� ���������	�B�-� f�Q���u��������� ����,P;` �q����������VERSI�@P�WQ d?isable^���SAVE ۅZ�	2670H7K69'�!4�0��po� 		(kR$�?;+2/ESeO/x/�/�/�/�*g,��/tz�n_�P 1ܸk�20
B�5<?N?��7�@URGE�B�P�^�aWFz0�QdT��pVW`�4LQ��W�RUP_DELA�Y ݼ��5R_?HOT %FnQ�3�O�5R_NORMAL�8�R
O_O.GSEMI>OdO�O�A_QSKIP3�p�+3x�O__0_ �M�5W_eWO_�_�_�_ o_�_�_�_oo'o�_ Ko9ooo�o�oYo�o�o �o�o�o�o5#E k}�U���� ���1��U�g�y���5�$RBTIF��4��RCVTMO�Uէå���D�CR3��I ���AC�}�C����C��?����>�9�<�<�Mä�`���2	1�$�,��� �(9���OC�?_ <
�6b<߈;����>u.�>*?��<���U���8?����� ��ߟ ���'�9�K�]�o���������ERDIO�_TYPE  �!=����EDPRO�T_CFG ��G�4BH3E����A2�� ���B� �T�b��� ��:�����п��c�� �O(�G_I�;�Y�[�m� �ϑ��ϵ������� ����E�3�i�Wߍ�{� �ߟ߱���	��-�/� ��?�e�S��w��� ���������+���O� =�s�a����������� �������K9o ]�������� �5#EGY� }�����/� 1//U/C/y/g/�/����/����INT �2��9J��ǱG;� ?&;s���N?�f�0 l?~;�/�? �/�?�?�?�?�?OO ,ORO@OvOdO�O�O�O �O�O�O�O_*__N_ <_r_`_�_�_�_�_�_ �_�_o&ooJo8ono \o~o�o�o�o�o�o���EFPOS1 1��̩  x �/:y�A?cN��x -?y����"� �F��C�|����;� ď_���������B� -�f����%���I��� �����,�ǟP�b� ���I�����ίi�� ������L��p�� ��/���ʿe�w���� ��6�ѿZ���~��{� ��O���s��ϗ� �2� �����z�eߞ�9��� ]��߁�����@��� d��߈��5�G���� �����*���N���K� �����C���g��� ������J5n	� -�Q���� 4�XjQ� ��q��/�/ T/�x//�/7/�/�/ m//�/??>?�/b? �/�?!?�?�?W?�?{? O�?(O:O�?�?!O�O mO�OAO�OeO�O�O�Ox$_�Cu2 1� �O�O_�_{_�_�O�_ s_�_�_�_2o�_Vo�_ zoo�o9oKo]o�o�o �o�o@�od�oa �5�Y�}�� ���`�K������ C�̏g�ɏ���&��� J��n�	��-�g�ȟ ��쟇����4�ϟ1� j����)���M�֯q� ����ϯ0��T��x� ���7���ҿm����� ϵ�>�ٿ���7Ϙ� �ϼ�W���{�ߟ�� :���^��ς�ߦ�A� S�eߟ� ���$��H� ��l��i��=���a� ����������h� S���'���K���o��� 
��.��R��v #5o���� �<�9r�1 �U�y���8/ #/\/��//�/?/�/ �/u/�/�/"?�/F?,_>T3 1�I_�/? ??�?�?�?�/O�?)O �?&O_O�?�OO�OBO �OfOxO�O�O%__I_ �Om__�_,_�_�_b_ �_�_o�_3o�_�_�_ ,o�oxo�oLo�opo�o �o�o/�oS�ow �6HZ���� �=��a��^���2� ��V�ߏz������ ��]�H������@�ɟ d�Ɵ����#���G�� k���*�d�ů��� �����1�̯.�g�� ��&���J�ӿn����� ̿-��Q��u�ϙ� 4ϖ���j��ώ�߲� ;�������4ߕ߀߹� T���x�����7��� [������>�P�b� ������!���E���i� �f���:���^����� ������eP� $�H�l���+�O�sY?k44 1�v? 2l� �/2/�V/�S/ �/'/�/K/�/o/�/�/ �/�/�/R?=?v??�? 5?�?Y?�?�?�?O�? <O�?`O�?OOYO�O �O�OyO_�O&_�O#_ \_�O�__�_?_�_c_ u_�_�_"ooFo�_jo o�o)o�o�o_o�o�o �o0�o�o�o)� u�I�m��� ,��P��t����3� E�W����ݏ���:� Տ^���[���/���S� ܟw� ���������Z� E�~����=�Ưa�ï ���� ���D�߯h�� �'�a�¿��濁�
� ��.�ɿ+�d�����#� ��G���k�}Ϗ���*� �N���r�ߖ�1ߓ� ��g��ߋ���8��� ����1��}��Q��� u������4���X����|������5 1�M�_���; A�_�����T �x�%��� j�>�b� ��!/�E/�i// �/(/:/L/�/�/�/? �//?�/S?�/P?�?$? �?H?�?l?�?�?�?�? �?OO:OsOO�O2O�O VO�O�O�O_�O9_�O ]_�O
__V_�_�_�_ v_�_�_#o�_ oYo�_ }oo�o<o�o`oro�o �o
C�og� &��\��	�� -����&���r��� F�Ϗj�󏎏��)�ď M��q����0�B�T� ���ڟ���7�ҟ[� ��X���,���P�ٯt� ����������W�B�{� ���:�ÿ^������� ϸ�A�ܿe� ��$� ^ϿϪ���~�ߢ�+� ��(�a��υ� ߩ�D�x�߳���6 1��� zߌ���D�/�h�nߌ� '��K�����
��� .���R������K��� ����k������� N��r�1�U gy��8�\ ��}�Q�u ��"/���/|/ g/�/;/�/_/�/�/�/ ?�/B?�/f??�?%? 7?I?�?�?�?O�?,O �?PO�?MO�O!O�OEO �OiO�O�O�O�O�OL_ 7_p__�_/_�_S_�_ �_�_o�_6o�_Zo�_ ooSo�o�o�oso�o �o �oV�oz �9�]o��� �@��d����#��� ��Y��}����*�ŏ ׏�#���o���C�̟ g�🋟�&���J�� n�	���-�?�Q���� ׯ���4�ϯX��U� ��)���M�ֿq�������7 1��ߧ��� �q�\ϕϛ���T��� x���߮�7���[��� ��,�>�x������� ��!��E���B�{�� ��:���^������ ��A�,�e� ���$��� H�����~���+�� O����H��� h���K� o
�.�Rdv �/�5/�Y/�}/ /z/�/N/�/r/�/�/ ?�/�/�/?y?d?�? 8?�?\?�?�?�?O�? ?O�?cO�?�O"O4OFO �O�O�O_�O)_�OM_ �OJ_�__�_B_�_f_ �_�_�_�_�_Io4omo o�o,o�oPo�o�o�o �o3�oW�o P���p��� ��S��w����6� ��Z�l�~�����=� ؏a����� �����V��ߟz����'���8 1�*�ԟ� ��� ��¯ȟ毁�
���� @�ۯd�����#���G� Y�k�����*�ſN� �r��oϨ�C���g� �ϋ�߯������n� Yߒ�-߶�Q���u��� ��4���X���|�� )�;�u��������� ��B���?�x����7� ��[����������> )b���!�E� �{�(�L� �E���e� �/�/H/�l// �/+/�/O/a/s/�/? �/2?�/V?�/z??w? �?K?�?o?�?�?O�? �?�?OvOaO�O5O�O YO�O}O�O_�O<_�O `_�O�__1_C_}_�_ �_o�_&o�_Jo�_Go �oo�o?o�oco�o�o �o�o�oF1j� )�M������0��T�:�L�MAS�K 1�W�N������x�XNO  �������MOTE�  ǌ  ��_?CFG ��O��l�PL_RAN�G ��q[��A�OW_ER �W�y��`�SM_DRYP�RG %W��%�����TART ��q���UME_�PRO�����H�_�EXEC_ENB�  �t\�GScPD��6�>�K�gTDBY�k�RMz��k�IA_OPTI3ONQ��^��INGVERS���Ȋ
�o�I_�AIRPURO� ���Մ1�m�MT_ Tl��`�OBOT_ISOLCŌ��-�4�0�o�NA�ME���n�OB?_CATEGňy��փ̀���سOR�D_NUM ?�q�*�H769  �t@�R��d�x�PC_TIMoEOUTQ� xx�oS232�1�ȅ�j� LTE�ACH PEND�AN���8����Ƽ ��pMai�ntenance_ Cons�r�����"���tNo Use�����@�R��d�v߈�v���NPO�ΐ��8�̥��C7H_L���^�J��	���!UD�1:1���R�VA3IL!�¥�\��_SR  �ʡ�8���R_INT7VAL���\��������V_DATA_GRP 2�ȅ��� D��P L�/�H�S�>�ȅv��� n��������������� ��F4jX�| ������0 TBdfx�� ����//*/P/ >/t/b/�/�/�/�/�/ �/�/??:?(?^?L? �?p?�?�?�?�?�? O �?$OO4O6OHO~OlO �O�O�O�O�O�O�O _�_D_́�$SAF�_DO_PULS����p[��SCA�N}���[���SC�m���`�Xj�
�p�p
��1�`��վQ�r H��_o o,o>oPo�_to�o�o��o�o�o����"ib2�d�Q�Qdx�a�
q�	�T�i @�7�FXjtv&y: ���t�_ @�sTʠ����~�T D��� +�=�O�a�s������� ��͏ߏ���'�9��K��߯�8wpZ�����n�  �ŏ;�o��ʑ��p�����
�t���Di_�jaѰ�X � �����U�Q 9�K�]�o��������� ɯۯ����#�5�G� Y�k�}�������ſ׿ �����1�C�U�g� yϋϝϯ���������	ߗ���2�D�V�h� zߌߞ߰�����e��  ��$�6�H�Z�l�~������}�0�r�� &�������)�;�M� _�q������������� ��%7I[m ������� !3EWi{� ������// //A/S/e/w/�ߛ/�/ �/�/�/�/??+?�� ����ibk?}?�?�?�? �?�?�?�?OO1O?I ROdOvO�O�O�O�O�O �O�O__*_<_N_`_ r_�_�_�_�_�_�_�_ oo&o8o,x�a�� Co�o�o�o�o�o�o�o �o"4FXj|���zmo���v���+����	�1234567�8]2h!BG!��%�\1}�k`�T�f�x������� ��ҏ��lo��1� C�U�g�y��������� ӟ���	��-�>��� a�s���������ͯ߯ ���'�9�K�]�o� ��@�R���ɿۿ��� �#�5�G�Y�k�}Ϗ� �ϳ����ϖ����� 1�C�U�g�yߋߝ߯� ��������	��-��� Q�c�u������� ������)�;�M�_� q���B���������� %7I[m �������� !3EWi{�� �����//// �S/e/w/�/�/�/�/ �/�/�/??+?=?O?a?s?�?McE��?�?�I/�?�?O�C�z  BpIj  � �H2_b } 6F�
[G�  	ĀAD�?�O�O�O�O�KDo�<�uO_$_6_H_ Z_l_~_�_�_�_�_�_ �_�_o o2oDoVoho �O�o�o�o�o�o�o�o 
.@Rdv� ������#��B��1iA�<� ��iA  ��/�I��v,�mAmAt  6@m����x�`�$SCR_G�RP 1�*�P30� �� ��A ��	 Ё�؂���1�����w��#��J�M��K@G�DCv����N�G��L	M�-10iA/8L� 1234567�890k@�� 8~k@MT20 ͐&-C
ș���A^H �؁Z�ǁ '�ǁ�C�G���-�	�v���������~ά��H�؀_�܇ǂ����5�G���o�A"����p�����^� h@_,V�l\@��B�%@�������9A6@ �  @�@8�L�N�?�^���H%@�q�K��F@ F�`�£Ϛ��ϲ��� ����!��E�0�i�� ��8�h�ߑߣߵ�B���X�	���-�� Q�<�N��r����� �����O�q�3�!�F��]@C�x��B`�8��>���~�6�i�@h8���%@���ȗ`�'��?-DA��H1a�]�> �A2��A T{��
ip���� (� � $��H3�l)J��Γ��ECL�VL  �A���7�?A��*S�YSTEM*�@V�9.10214 ��8/21/20��A �@�z��SERVENT�_T   $ �$S_NAME� !	 POR�T�@!ROTOz! �_SPD  ���/ TRQ   
,#/AXIS5!:'2 � 2c�,#DET�AIL_  �l $DATE�TI! ERR_�COD�#IMP_wVEL4@ 	�"�TOQ�$ANGL;ES�$DIS��&�" G%%$LIN��" +$REC5!� ,!O%i � M�RA�! 2 ]d2IDX!�$�B  �0$O�VER_LIMI� I 	��,#OC�CUR5!  ��+COUNTE�R�%FZN_CF�G5! 4 $�ENABL�#ST�� "FLAG"D�EBU�3R�! �ѐ~3��5! � �
$MIN_OV;RD�@$I�� x�2�1�5FACEe"��1SAF�7MIX�EDL�9�!�2RO�B%$NE&AP�P�"�SHELL��4	 5$�J?@BAS�#RS�R_�5  $�NUM_y@�  �xA1�'y@2�J3��J4�J5�J6�J7r�J8�'lAROO �� CO�ONLY��$USE_A�B#xBACKE�NB�  PIN>0T�_CHKSOP_�SEL_�0,Y_P�U;Qo1M_�!OU#PNS|F PYC�&��0EPM�%TPFWD_KAR�! P�!�RE$$OPT�ION�2$QUEԃY" D�RYRB$C�STOPI_AL;SYCEX+STQ�P�$[XTSPM1i2"�MA�1STY;TSmO
`NBRDIGQ�TRI�3�Q�WIN�I�M& 8bNRQ�xf`ENDNd$�KEYSWITCaH�S�QZa�THE�P�BEATM�SPE�RM_LE�"�QE�� �gU�SFd�RS~_dDO_HOM�09ORA/PEFP !"0L�3U ST�bRC�`�OM�#�!OV_M�SJQ ET_IOGCMN+S�W5a��XEHK !
 D ��7qSU�"�RM�P+S� PO7B$�FORC�SWAR�Nk|OMrP ~7�$FUNC�2�3U	0}QAR'`�u�2�v3�v4�q�W��SC0O�PL�ry�"�XUNLOeP��$:�ED� ���SNPX_AS�2 0�@ADD|�0�1$SIZ�!�$VAR�'MU/LTIPRZ��p�A�q � 1$tY[�r	�B`��"�AC� ΆFRI	F">0S�P�y"t���NF{dODBUS_ADw2�B��&�CM�aDIA�q$DUMMY15ajM�3J�4J��Sz@>  � x��"�TEqM�8J�SG�L��TAJp  &�0���@J������STMT�Q��PS3EGb��BW�P���SHOW��!BA=N̐TPOF�M��9J�0J�(a��SVC�G�2 ��$PCpP?0-�G3�$FB�qPD�SPb�PAFPF�L VD/�~�2� ��!A0��@� ���p��@�p��	������5��U6��7��8��9��A��B���p��h ��Ր��F���P���T��P���l�P�̩1٩1��1�1 �1�1��1'�14�1A�1PN��!ǘ�2��2��U2��2̩2٩2�U2�2 �2�2�U2'�24�2A�2N�U3��3��3��3��U3��3̩3٩3�U3�3 �3�3�U3'�34�3A�3N�U4��4��4��4��U4��4̩4٩4�U4�4 �4�4�U4'�44�4A�4N�U5��5��5��5��U5��5̩5٩5�U5�5 �5�5�U5'�54�5A�5N�U6��6��6��6��U6��6̩6٩6�U6�6 �6�6�U6'�64�6A�6N�U7��7��7��7��U7��7̩7٩7��U7�7 �7�7�U7'�74�7A�7N���"VP�`U3"# < �B
�� ! x $T�OR�Q@�  �"Mb$ R1 L@BQ_W0AR��%T!�p�$S[iC�Qp�_U����rYSL�   � x���7���m��0���`�R�VA�LU�5QP�V]�F��ID_L�"%H�I*I�r$FILcE_xSM$BD$s��SA21 h�5y E_BLCK��S�"���(D_CPU�)y��)m��3P/b$�Y�Y��rSR ? � PWY0Pl�� 1LAƑS11�314RUN_FLG(54,14�`/5M14M15HrP4o0�4��T2�Q_LI��r  k@G�_Ob�PP_E3DI+RT2 @�3�20�$P�!������TBC2x� �}�8P/0T�QƏ1FT'dD5cTDEC/0A`a�0@M	��F.AGTH����DDOPGRQH��pERVE(crD5crDa���14PG@ �X -$�ALEN`(c�D5c�@`RA�PLF��W_k�#1�A�:$2�GMO�!C�S�DPIZP�F!Y8̝@![DE1U�LA3CEXrfCCB���`_MA^�0VjU@W�jQTCVq\�Q@WT �a�Z�U�Zd�/S]��UT@S]�J@`AY�M�T" Jjgv�/Ua@U�A2)pp\�5a.S6H�JKHfVK$�ZaU�Zaa�O`J�ra^c�JJfcJJncAAL^c�`fc�`�fm��b5OC�PN1�\�`�[�nP�L
P_�� �� �1CFb� =`5GROU ����P�N�0C�� pR�EQUIR]B�E�BU̓�A�V$T1P2Vq�@@v�1a���4 \�p�8AP�PRLpCL�
$:�0N�xCLO�0�y�S:E�y/U
�1�� ��0M,@oP�PF�N�t_MGI��pCx��z �d�lP�BRK��NOLD��R�TMO�1I�6��uJ�0H�P�dLPfcLPnc�LP�cLP�cLP6��7ă���;`�B�4G� Ir�B$��<U��PATH��@����H��p[p�.�SCA�2L��r�qIN�BUCP�A\�-Cf�UMe�Y�@� `l�&!xA�����������PAYLOA�D�J2LR_A	N$AȓL0ҙΑ�ޑ�R_F2LS3HRlD�LOӔ[���i��i�ACRL�_�!Y�L�U���gbH���$H�z�F�LEX�s�0BJ�6 P�r�?
OqO��Om"���E  :�O�F@P�#��O�a0@P�O�O�LF1#�q� ���O__0_B_T_��E^_p_�_�_�_�_�_ �_�_�ȩ��WcHd��@��o!o3o"�:jT����XraFe���Qe Z�3�]ooo�o�`�e�e��e�e�o�o�o�i�1BJt! ��0#5 AT��Hq�PCEL�T1p�OxJ[p� VpJE3�CTR�U���TN)l�@wH�AND_VB���� ׄ" $��Fi2�<D�SW�g��v#� $$M ��yM#��2�-�O� �q�K�A) ���v(!Dh� �A��#�A1�AA@�s��� #�D1��D@�P �G"0		S�T%�2�NC�DY.0�p�T�{����@ �#�����Hg��K�-�G�P����������ฅ��ʂ��5$ ���� Ʊ�q�ASYM0���Ip0�#wL��P�_ n0A�a�t�^�`��~�������ƓJ͜~�ߚp������_VI���<(�sM V_UN �2; b#��
�JIez" �z"�~$4��$�&=���PP�~�_�q�5;�|�������T�03HR�0�1%��01L���2DI@�;sOO4q �110�& ��
��IeA��4�|1�����3��|�0�20 �' � ��M�E���Х2�"�TC0PT����1�`��d����8�1�9T���a $DU�MMY1��$P�S_��RF^�`0u$(F�pFLAp�YP2�BB�3$GLB_T�E5]E�0ౡ��۰��1( XX�p@wׁST��Vp�SBR�M21_�V bT$SV_E�R�O��C�CCL�w@�BA�O2,0G�LD EWq) 4\p�1$Y��Z��!WS>`���A�0e�t`2�AU�E* ��yN P�$GI��7}$�A �@�CPq+ LpAV��}$F�EIVNE+AR�N��F�Y��TANC��  ��JOGR�t� �,�$JOIN�T=�N��a�AMSE]Tq-  >WEvU�:�SA�+1^Q;�q_.� ��U���?�VpLOCK_�FO���K0BGL�V��GL:hTES�T_XM�p�QEM�P�P��^buB%`c$U��B=�2*Vp�S�a+Ob��*`�a)ƥACE�`RS�` $�KARP�MQ3TP�DRA�@�d�QVE�C4��f�PIU�a,��aHE,`TOOL�e��cVd�RE�`I�S3�r6����ASCH�P[p-qO>���3D3��QPSI��r  @$RAIL_BOXE=ѽ�@ROBOUd?���AHOWWAR���tq%@@qROLM 0B�u �=t�r0�bp��nـO_F1�!�@�HTML5D1U����@2qځ/�^*0R
�`O��0�R]��Q�p�)VOU�R1 d��@�e)�v�P�%`/$PIPVfN0�r�br2q���a�p�CORDED*`6���P�XTV�DQ),0,�O��0 2 D \@OB��z�*`�����C[@���|�SYS���ADR{�,0�0T�CH:� 3 ,���EN52��A1a_�AT�	��,0V�WVA�14 �� �`�BE5PRE�V_RT�$E�DITT�VSHW�R1��Fs�� Q�< D�0�����$HEAD�� ����\�KE Q@C�PSPD��JMP���LD5��R�g4Q5�����I_`S{�C��NEp|��T'ICKe�oM�����HN�A6 @p����Ñ_GPR��Yv��STY	�>qL�OwA�B�N� �7� t 
O�G�%�$4�AT=�@Sq�!$p!=м1HEy0GF9PRR�SQU�`X�<IB;!TERC�0��z�S�8 HP��@.�0�-���a^�O�0�3��IZJDAQFE$APR��1Ap����.�PUAဵ_DO��R�XS�PKD6A�XI���s�aUR I��|�{p@�͆��J�Y_�`߂ET�P3b���5��F5��A,B8D9Hw���Up�SR��9l ��M�%�[�8�m� K�[�V�[�d�[�t��� ���Ŧ��Ŷ������������!��C6���C��ͯ����ASS}C_@ : h�@cDS`��a@SPv0&��AT��L���?���BADDRESzsB_�SHIFA�^{`_2CH{�Ɂ�I~@��TU~@I�*� ;�RCUSSTO��VbIj2A< �Gh��d�
^j�
��V-����0= 	\�@G����o�>�����C��A��~�F��B����TXSCRE�E��><0��TICNA�COP��AT,�8���? T���@ d�߁�A�@L���ނ��H�[�RRO �Pހ���E�5{@UE�@# �M��6@S�A߁'RSM?���U��
�D6��00S_S��i ������i�Cb���3� 2?��UE�Ap2�Bp�GM�T� L�!���@O~�U�BBL_Bp9W�0�0B ���v5OQ�LE�xzpE�RIGH��BRD�D�CKG�R�0�T����WIDTHHs��ĲUq|BAq�UI�pEY�Щ1C6��p�p�bpl�BACKЀ�0B1�A�0FO��DLAB��?(�0I@p#b$URL�qqCO	�0Hl� D 81�P_����0R P%b/ÐHx Aa0�O�0E�I��G� U� �R3b�qLUM�Ķ�GERVM��@
P�PjF�0�GEu0{Q������LP4%
�	E���)Q'��_(�Ѩ_(,p^)5\+6\+7\+8A"��3k��P���F,qaS��E�	USR�DG �<�@�0UERT�ERF�OB�ERPRI�mxLp�!30TRIP^qm�UNDOg5H<PàL0���qڗ8{bްؠ I�� .o�G ��T�p��L �2OS�1�6R�r�v3�a�AJ�OS^��2b��u4U<!�AK��?�?��<"a�v3OF�FT`�@L�@�3OU@ 1J�@?DgD-K�@GUفPfA�Rp�C}ьGSUBb���@/ SRT�0B�M0I��Q�pO�ORBp�E'RAUT��DT�I�r�A_R��N |]���OWNy0�$GSRC}�����DT`<>UR�MPFIy�y��ESP|�G��u #��'rLARm�67O `@WO����=��COP!A	$հ{0_YPr�Q.��UWA_�Cra�Q�P��S�Qr&�4��rW� �P?�SHADO�W��s"a_UNS�CA�c"c�/cDGyD7q��EGAC�Sld�'�PG�Q�N��STE���O���t�PE"��VuWDt�TRG��6R �>��jMO�VE}�#A�bANG����f-C�f�3�bLIM_X!Cv'Cv�h q|��g?06��`"B�VF���C��VCCԢ��S?�C��RAध�`ϥD��@NFA��R@�]�E,�Q2>0G����R:�{0DE�b
�p���p6T� i�؁ϣA�u�㡹W C% ��DRI�`��aV�[�*��S�D�$MY_UBY�$�}�3ϥ~������Q���P_8`y���L��B�M�$�DEY�
�EXc ���UMUbِX�d����US��˰.0_R�"B#06�z�fG�PACIqt �`HQ�dI�-CI��3I����QRE���1�Bq�sI��U ?�
�PG�`P�⎐G0�s	R�0�V�k��ҲB	�R��R�dSWHA�os�@��n�O�!��A��[�E� Uȑ��a�@�0�sHK
��W���aS���Q��cEANS��P�x�@�rMRCV6WX �- O�pM��C��	��?C����REFb������
r� ِ0��ꡨ�꡹����A�_;PW�B�o��� �`��k�\���x�Q�r3Y ��a��ϒ��1`�$GROU@���3��¶�s�pT��
��20$ ����0X �V�Ӂ�ֱ���U�L�qW�PC%p�X��NT�S+ĔR@*��6��!6���L��@_Ű�_��k��!�p�TIЙ�Z t@M}D�@AP_HUx���`��SA�cCMPB}�F�����Ų�_��ARqty���W�j�X����VGF`S[� �M0����UF_{�˂��@JʼRO� T�շ����|.�URE9��6�RI;���I&༨�o��o{FQyFQ'C`wIEN�H��xx� V�1 ,r��A��?�W�|���Q/��V큂��LO�p'�\ax �����!N{SI"VIA_�R�;�\ �� HDR{ )$JO� �b�$Z_U�P)p��Z_LOW �������\(p���P鱬3�9���Ⴐ���'Q�����"�]o� 0�PA�{ �CACH�� ��}���퀙�!�P]S�C(qIB�F#���T8� ��|�$HO�1R��/�%�"f�������?�RQ0!��cPVPx��� H_SIZ�RZ��M��N�Q�sMPr
�qIMG�d���AD�	�RMRqE���WGPM�p�NDRP�VASYN�BUF�VVRTD�� W��OLE_C2D,tc�1@C�q�Uۃ��Q��EC;CU{�VEMe�}�<d��VIRC�0�
" {�LA��RQX}0\0��AGR�GXYZ)��C�W�� �����A�T�p܂�IM��G`��G/RABB�1Y�b��� ���^q`
�CKLAS��b�Y@'_  񱵵T��5P�@�21T$b��p!�`� ���SP�G�%T@Q�RQ�q�P�"x�I�$�|��=�BG_LE3VE�QL�PKL��l"ѥ�GI� NO�Q�q2,�͐HObPRa � �F����bE6S��g]2RO�cACCEe@����x4VR�A�y1܂R`6� AR�cPA@�>���D�SREM_B�Q$ ��͐JMP�U�XAbi$1�$SSlSFD ��p͐��|�Y@c  ���S� ��N/D`LEX�&dbSdqg`��&DR�w$YQqH(`hqH҄�cABP2h��e� �є`V|��cPMV_PI���DX�`�@3����IF&�\rZ�JT�E�@��0�H���E�AGAU?��LOO�d?�JCB�TZ�'B`H +cPLCAN'r��L2��Fw ��D?V5Y �WM��~Ppu�T�FS��U�Q �ѥU����V2DbX9�1LRKEZq�1�VANC]C�R_9O�|`f (�p8��s$\�3Zr�rR_}A3� g 4���dovn#p� �_���h� h��9��ĬvOFF�sfW@������EA��
� LSK���MN��q�g �S`��|@c"i < �WJ��=�UMMY�Y���n�D�P��}�CU��1�U��pj $�TI}TV1$PR8Af��OP����SF����Cki �|6���.�!SMO!�l%BXCb�4J�p��ZD�vgm DQx�AL^1#IM; ��0IN�_MSG_Q�SHwЅ_pn%B­w8�%�M� �X�VR"�oI"�pT��5 �ZABC���p��Ƃ��Ӡ
�AA%��`VS.� q � w0���=�CTIVeAI�O�b�	s�ITVlLW�DV@
l�"��2� DI�� @�� ��|A��d���N�LSTs���ݰ��7_ST��Pa%��DCSCH��r LQp�����~P1��m�W GN����r���_FUN�� ��7ZIP!�s%B� �L8�L|�Ѣu�Z/MPCFʅt�r9����L�DMY_L�N$pq
8�'�˄u $��Q��CMCM��CLCOART_����P�a? $J����D=��¢��u�ǥu����_�p���U�X�P�UXEUL ����
�̥
��.�8�>���FTF����k�����Z�v� �*�@��Y�%�D.  w 8/ $R� U�Q���EIGHe3�x?(��0��0��p��A$x� �=0�sq�$B������b_SH�IFB�	�RV�PFL��1�	$)0C�� �����d�pl��r�"�l��D|ȕ�C �N1V�a���PH�0%чy ,�0��ֿ� ��$S{0DEFA�Un�t�����������HO�T������MI�POWERFL �Oa����%�WFDO�� ����Y�~�`1 ���qѾ� L!ip_�EIP5ԑ����j!AF���`�߼�O!FT������f�!��-����.S�!R9MHQp�7�B��f�@o�5�������!OPC3UA�����7�!TPP�@8���yd&���!
PM�p&�pXY����er����J����f��!�RDM-@V��g|
g!R90h2��hV�!
h�~������i��!R�LSYNC &�8�K!ROS̉�r�4:�!
CEL�MT�`��֙k��!	��PSd���l�//!��WASRC6��m�/{/!�USB�|/��nj/�/!S#TMP��/��o�/?@�7?*?`=e�I���KL ?%q� �(%SVCPR#G1`?�:�52�?�?"�03�?�?�04�?�?"�05 O%O�06HOMO"�07pOuO�08�O�O�09�O�K�4~�O �1�?_�1�?=_�1�? e_�1O�_�1:O�_�1 bO�_�1�Oo�1�O-o �1�OUo�1_}o�1+_ �o�1S_�o�1{_�o�1 �_�1�_E�1�_m �1o��1Co��1ko ��1�oe?w2�0~?�0 0�u��1y��������� �Џ	��-�?�*�c� N���r�����ϟ��� ��)��M�8�q�\� ������˯���گ� ��7�"�I�m�X���|� ����ٿĿ�����3� �W�B�{�fϟϊϱ��������k:_DEV� q��M{C:�4���?GRP 2q�����0bx 	�/ 
 ,c��|� <�hߥߌ��߰����� ��#�
�G�Y�@�}�d� ����������d� 1���U�g�N���r��� ��������	��? &cJ����� ����;M4 qX������ /�%//I/0/B// ��/�/�/�/�/�/�/ �/3??W?>?{?�?t? �?�?�?�?�?O�?/O AO�/eOO�O�O�O�O �O�O�O�O_ _=_$_ 6_s_Z_�_~_�_�_�_ �_HO�_'o�_Ko2ooo �oho�o�o�o�o�o�o �o#5Y@}d v�
o����� 1��*�g�N���r��� �����̏	���?� &�c�u����P���ϟ ���ڟ�)��M�4� q�X�j�����˯��� ��%�|��[��� f�������ٿ����� ��3��W�i�Pύ�t��ϘϪ���7�d ���	���	�B�-�f�Qߊߙ�%��߾�>�����у����� ������9�'�]�k� �ߐ���S������� �����;�}�b���+� ��������������C� i�:y�m[� ��� ?�3 �CiW�{�� ��/�///?/ e/S/�/��/�y/�/ �/?�/+??;?a?�/ �?�/Q?�?�?�?�?O �?'Oi?NO`OO9OO �O�O�O�O�O�OAO&_ eO�OY_G_i_k_}_�_ �_�__�_=_�_1oo UoCoeogoyo�o�_�o o�o	�o-Q? a�o�o��o��� ��)��M��t�� =���9���ݏˏ�� %�g�L�����m��� ����ٟǟ��?�$�c� �W�E�{�i������� կ���;�ů/��S� A�w�e���ݯ¿Կ�� ������+��O�=�s� ����ٿc��ϻ����� ��'��Kߍ�r߱�;� �ߓ��߷�������#� e�J���}�k��� �����+�Q�"�a��� U�C�y�g�������� ��'�����+Q? uc�������� �'M;q� ��a����/ /#/I/�p/�9/�/ �/�/�/�/�/?Q/6? H?�/!?�/i?�?�?�? �?�?)?OM?�?AO/O QOSOeO�O�O�OO�O %O�O__=_+_M_O_ a_�_�O�_�O�_�_�_ oo9o'oIo�_�_�o �_oo�o�o�o�o�o 5wo\�o%�!� �����O4�s �g�U���y������� �'��K�Տ?�-�c� Q���u��������#� ����;�)�_�M��� ş����s���o�ݯ� �7�%�[�������K� ����ſǿٿ���3� u�Zϙ�#ύ�{ϱϟ� �������M�2�q��� e�S߉�w߭ߛ߽�� 9�
�I���=�+�a�O� ��s��������� ���9�'�]�K����� ����q��������� 5#Y�����I� �����1s X�!�y��� ��9/0/�	/� Q/�/u/�/�/�//�/ 5/�/)??9?;?M?�? q?�?�/�??�?O�? %OO5O7OIOO�?�O �?oO�O�O�O�O!__ 1_�O�O~_�OW_�_�_ �_�_�_�_o__Do�_ owo	o�o�o�o�o�o �o7o[o�oO=s a�����3 �'��K�9�o�]�� ���̏������#� �G�5�k�������[� }�W�ş�����C� ��j���3��������� ������]�B���� u�c������������ 5��Y��M�;�q�_� �σϥ���!���1��� %��I�7�m�[ߑ��� ���ρ���}���!�� E�3�i�ߐ���Y��� ����������A��� h���1����������� ����[�@�	s a�����! ���9o]� �����/� !/#/5/k/Y/�/��/ �/�/�/?�/?? 1?g?�/�?�/W?�?�? �?�?	O�?Oo?�?fO �??O�O�O�O�O�O�O _GO,_kO�O__�Oo_ �_�_�_�_�__oC_ �_7o%o[oIoko�oo �o�_�oo�o�o3 !WEg��o��o }����/��S� �z���C�e�?���� я���+�m�R���� ��s�������ߟ͟� E�*�i��]�K���o� ������ۯ��A�˯ 5�#�Y�G�}�k���� 	�ڿ������1�� U�C�yϻ���߿i��� e���	���-��Qߓ� x߷�A߫ߙ��߽��� ���)�k�P���� q���������C� (�g���[�I��m��� ����	��� ������ !WE{i���� ���	S Aw���g�� ��///O/�v/ �?/�/�/�/�/�/�/ ?W/}/N?�/'?�?o? �?�?�?�?�?/?OS? �?GO�?WO}OkO�O�O �OO�O+O�O__C_ 1_S_y_g_�_�O�__ �_�_�_o	o?o-oOo uo�_�o�_eo�o�o�o �o;}obt+ M'������ U:�y�m�[�}�� ��Ǐ���-��Q�ۏ E�3�i�W�y�{���ß ��)�����A�/� e�S�u�˟�¯��� �����=�+�a��� ��ǯQ���M�˿�߿ ��9�{�`ϟ�)ϓ� �Ϸϥ��������S� 8�w��k�Yߏ�}߳� ������+��O���C� 1�g�U��y������ ������	�?�-�c��Q�����������$�SERV_MAI�L  �����~��OUTPUT��_��@���RV 2w�  �� (��I���SAVE��TO�P10 2#	 d ���� ��'9K] o������� �/#/5/G/Y/k/}/ �/�/�/�/�/�/�/? ?1?C?U?g?y?�?�?�w�{YPf��FZ�N_CFG w���W~�1GRP 2�7�t ,B   �A'@��D;� B}(@�  B4��RB21VH7ELL�2	w�r�6 7�7�O�K%RSR�O�O�O�O�O _�O3__W_B_T_�_ x_�_�_�_�_�_on?�  ��Ro�Ko]o+bio ���eo�b�`�bg3b2���dultm�bRFHKw 1
`K �o 0YTfx ���������1�,�>�P�LLOMM� `O��QBFT?OV_ENB��+�r�bOW_REG�_UI����IMI_OFWDL�����*E��WAIT�� �i�2����*�wTIM���T��VA��+���_UNcIT����r	LCڀWTRY�r���MON_ALIA�S ?e��2 he���!�3�E�S��� v�������W�Я��� ��ï<�N�`�r��� /�����̿޿𿛿� &�8�J���[πϒϤ� ��a��������"��� F�X�j�|ߎ�9߲��� �����ߥ��0�B�T� ��x������k��� ����,���P�b�t� ����C����������� (:L^	�� ���u� $ 6�Zl~��M ����� /2/D/ V/h//�/�/�/�/�/ /�/
??.?@?�/d? v?�?�?E?�?�?�?�? O�?*O<ONO`OrOO �O�O�O�O�O�O__ &_8_J_�On_�_�_�_ O_�_�_�_�_o�_4o FoXojo|o'o�o�o�o �o�o�o0B�o Sx���Y�� ����>�P�b�t� ��1�����Ώ��򏝏 �(�:�L���p����� ����c�ܟ� ��$��Γ�$SMON_�DEFPROG �&���N�� &*S?YSTEM*+�o�����?=�R�ECALL ?}�N� ( �}!�xyzrate �124=>169�.254.��12�0:19636 ���ɠȡ�����}
��1 ��ǯٯj� |���!���;���_�� ��'�ο˿ݿnπ� �ϥ�L�I�[������ #ϵ�����j�|ߎߡ� ��E�W�������1� ����f�x��߯�A� S�������-���� ��t������=���a� ����)���8��p ����NK]�  %���l~� �5GY��/!�:copy fr�s:orderf�il.dat v�irt:\tmpback\��d/�v/�/1*"mdb�:*.*?/Q/6 `\/�/�/?$5x*$:\�/40�/��/q?,�?�?}6*5a2?D? ��?�?O/1/�/U/ fOxO�O�/�/JO�/�O �O_?-?�?Q?�Ot_ �_�?�?<_N_a_�_o
�_� �_�_�_ko�}o�o��17572�]o�o %�o��o�ol~�#Imd�:picksim�_part1.tp�Eemp�OFs� ���o�o?z��o������&ptpdisc 0N�GrI�[������#stpc?onn 0 Ϗŏ�׏h�z���w2�uomay�P�Ip]�� ����2��ɟ۟l�~���#�d��E�W�� �������6�ȯگk� }���"O4O�OX���� ϠO�OͿFsܿm�� ��$_7oIoC�a����0�ϩ_����2 ��r� ��ߩ���D�_���� �'���K���n�����p�$SNPX_�ASG 2�������o  0�q%������  ?���PA�RAM ����� �	��Pʠt�p��1������OFT_K�B_CFG  ��s���OPIN_�SIM  ���,����������R�VNORDY_DOO  6�b����QSTP_DSB�v�,���SR ��� � &�0�Q�w�tG�TO�P_ON_ERR�����|PTN ���� �A��RING_PR�M���VCNT_OGP 2x�.���x 	
	�p�0�T��VD� RP' 1�/�E�� 7������� //1/C/U/g/y/�/ �/�/�/�/�/�/	?? -???Q?c?�?�?�?�? �?�?�?�?OO)OPO MO_OqO�O�O�O�O�O �O�O__%_7_I_[_ m__�_�_�_�_�_�_ �_o!o3oEoWoio{o �o�o�o�o�o�o�o /Ahew�� ������.�+� =�O�a�s��������� ͏����'�9�K� ]�o���������ɟ۟ ����#�5�G�Y��� }�������ůׯ��� ��F�C�U�g�y��� ������ӿ��	���-�?�Q�c�mPRG�_COUNTW�9���ENB����M��Y���_UPD� 14T  
xϣ���/�X�S� e�wߠߛ߭߿����� ���0�+�=�O�x�s� ������������ �'�P�K�]�o����� ������������(# 5Gpk}��� �� �HC Ug������ �� //-/?/h/c/ u/�/�/�/�/�/�/�/ ??@?;?M?_?�?�? �?�?�?�?�?�?OO %O7O`O[OmOO�O�O��O��_INFO {1����P	 �O__@_�+Y@l�@Iʟl?Z�F_-S��̵��5A�u�9	�]�Ǝ�@�K]�A���@CP A!" ?�nn_��A D5Oy����C����($6�T�5+���Q� �8�h�Ca���.~:��1�５���YS�DEBUG�������@d��
`SP_PwASS��B?k�LOG �F.�  �@�X�O�  ����AU�D1:\Hd�NIb_MPCNm���o�o����a�o ���fSAV Qi��2Qqal�b�E�hSV�k�TEM_TIME� 1Qg� 0o`2T��Z����^sMEMBK  	����q`qo��� �X|��� @ ��C�"�G�W���z�����a 2[@}q��я���/s���1�C�U�g�y� �{�����ß՟�����/�i�e>�c�u� ��������ϯ��� �)�;�M�_�q���������\uSK�p�x��`������.�@e���2,�W�AW�A�9t��i��Ϧ�(��#!������� ���<�-�� �-���0`F�t߆ߘߌ�Y΀��������(��@$,�P�D�t��� �����������(� :�L�^�p��������������T1SVGU�NSPD2e '�e���2MODE?_LIM �vvqd b��2��Qm���ASK_OPTGION`�y aS�_DI+`ENB � b�esBC2_GRP 2ܵ c|r�[R��C������BCCFG �7| (��b�L_U@R� v������/ -//Q/</u/`/�/�/ �/�/�/�/�/??;? &?_?J?�?�?7ց<�? �?�?�?p?�?+OOOO :OsO~�O�th@�O�O �O�O�O	_�O-__=_ ?_Q_�_u_�_�_�_�_ �_�_o)ooMo;oqo _o�o�o�o�o�o�o�h �03EW�o{ i������� ��A�/�e�S�u�w� �������я���+� �;�a�O���s����� ͟��ݟߟ�'��K� c�u�������5�ۯ ɯ����5�G�Y�'� }�k�����ſ��տ׿ ���C�1�g�Uϋ� yϛ��ϯ�����	��� -��=�?�Q߇�u߫� a����������;� )�K�q�_����� �������%��5�7� I��m����������� ����!E3iW �{����� ��#5Sew�� �����//� =/+/a/O/�/s/�/�/ �/�/�/?�/'??K? 9?[?�?o?�?�?�?�? �?�?�?�?OGO5OkO !�O�O�O�O�OUO�O �O_1__U_g_y_G_ �_�_�_�_�_�_�_�_ 	o?o-ocoQo�ouo�o �o�o�o�o�o) M;]_q��� �O���%�7��[� I�k������Ǐُ�� ���!��E�3�U�W� i�����ß���՟� ���A�/�e�S���w� ��������ѯ���+� �C�U�s�����������˿�߿���3���$TBCSG_G�RP 2���  �3�� 
 ?�   ^�p�Zϔ�~ϸϢϴ�@�����$�7�>�E̿d0 �S�?�3�	 HCA��"�>l�"�CS�BpVߙ�c�u߇����B�$�>������"�Bl����)�A������G�"�;�B�)�+�Q�G��$_��A3�"�Q���T��Ѩ��@����� '�:���e���M�_�x������?�ff��� ��	V3.0}0V�	mt2 * 2�$��<23�G�� [ -\  q��7�+J2>�E����CFG !��eO� R��
����0� 0Vd�d�u� �����/// P/;/t/_/�/�/�/�/ �/�/�/??:?%?^? I?�?m??�?�?�?�?  OOV�p�O/OAO�? tO_O�O�O�O�O�O�O �O_(_:_L__p_[_ �__�_�_3���_�� �_ooIo7omo[o�o o�o�o�o�o�o�o 3!WEgi{� �������-� S�A�w�e�����m�ŏ ׏������=�+�a� O���s�����͟ߟ�� ���9�'�]�o��� ��M�����ۯɯ�� ��5�#�Y�G�}�k��� ����׿ſ����� C�1�S�U�gϝϋ��� ������	����?�� W�i�{�%߫ߙ߻߽� �����)��M�_�q� ��A��������� �%���5�[�I��m� ��������������! E3iW�{� �����/ ?AS�w��� ����/��O/=/ s/a/�/�/�/�/�/�/ ??�/%?K?9?o?]? �?�?�?�?�?�?�?O �?!OGO5OkOYO�O}O �O�O�O�O�O_�O1_ _U_C_y_g_�_�_�_ �_�_�_�_o	o+o-o ?ouo��o�o�o[o�o �o�o;)_M ����w��� ��7�I�[��'��� �����ُǏ���� 3�!�W�E�{�i����� ����ß�����A� /�e�S�u��������� �ѯ���o1�C��o ����s�����Ϳ��ݿ ��'�9�K�	�ρ� oϥϓ��������Ϲ� #��3�5�G�}�kߡ� ���߳��������� C�1�g�U��y��� ������	���-��Q� ?�a���u���%�W��� ������M;q _������� #%7m� �]����/� /!/3/i/W/�/{/�/ �/�/�/�/?�//?? S?A?w?e?�?�?�?�? �?�?�?OO=OOO�� gOyO�O5O�O�O�O�O �O�O_9_'_]_o_�_ �_Q_�_�_�_�_�_�^�  %`)c �)f=o)b�$TBJ�OP_GRP 2�"�U� _ ?�)f	Ub�\c$cl��P��pJ�`��xe  � �� � ��`�)d� @%`tb	 ��CA��f��S�C��_)eta�b3�33�f�oz=�_��CS�?��Y�1ru`B�;pp�gLWw�o�o?�a�u�ޜz<؄-r��a��u=�)eB��w?C�  D�a�o�#�-�;��B9l�`2u�ff�n�&)eAЇ��w���>��ͭ�����;�ǎ���@fff���b�]���A���������9�ˌ�X��@�o�폎������%��ɟۛ;������@�o��� {����9�1�g�Y�C� Q������E�ϯ�ӯ ��@��կ_�y�c�Pq���пct�)f���	V3.00�zcmt2��*��yd$a)�4� �F� G9| �G�v�G�/��G�� H�@�H,�H.���HC� HYA@�Hn��H�� �H�� H�Y@�H�`H����H�c�H��H̿�H�nD��G G.A �GKm Gh� �G��G�x��G��G����G�:�G�Ѐ�G�f�G����G��\��H
�_�H��H���H @�H'��d�ր=L��=#�
������)bQ3o�+�)f/��?�߀f�d�RcESTPARS�hn`�RcHR��ABLEW 1%ci�)d�_�D� �@$�_�B_�_�(g0a_�	_�E
_�_ؾ�)a_��_�_�����RD	I��ma�����������O������������S��kc  I���������� *<N`r��� ����Hm���� lb��C,�>�P�b�� �2�D�V�h��)N�UM  �U*ma�`1` ������_CFG &�+��a@U`IMEBF_TT�Ѻkc��T&VER�Uj&�T#R 1'��' 8&�)b$`�! �PN  �/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? <OO)OrOMO_OuO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_4oo!ojo EoWomo{o�o�o�o�o�җ!_!�&@�%���MI_CHAN�`' �% .sDBGLVL`'�%��1p�ETHERAD �?���p�/���o�o��y�1pRO�UT~ !�!��t��|SNMAS�Kyx�#�q255.?��=�O�a�Á��OOLOFS_D�I���ecyORQCTRL (�+��0�ߍTΏ��'� 9�K�]�o��������� ɟ۟����#�3�͏�V�E�z�~�PE_D�ETAIWx��PG�L_CONFIG� .)"!���/cell/$C�ID$/grp1�~�����*�<��� �g�y���������P� ���	��-�?�οc� uχϙϫϽ�L�^��� ��)�;�M���q߃� �ߧ߹���Z����� %�7�I��������������M}n��!� 3�E�W�i��k���p��m���������  g�DVhz��- ����
.� Rdv���;� ��//*/�N/`/ r/�/�/�/�/I/�/�/ ??&?8?�/\?n?�? �?�?�?E?�?�?�?O "O4OFO�?jO|O�O�O �O�OSO�O�O__0_ B_�Of_x_�_�_�_�_��_͠�User View ��}}1234567890oo'o9o�Ko]oed�`£�o���Y2�Yb_�o�o�o�o !�o�o�R3�oo �����(��n4^#�5�G�Y�k�}�����n5�׏���@��1���R��n6Ə ��������ӟ�D���n7z�?�Q�c�u����������n8.�����)�;�M���n�t� �lCamera�Z꯳�ſ׿������E��7�I� [�ouχϙϫϽ���ŉ  ���i���1� C�U�g�y� ϝ߯��� �����	��-�?�f����]y�ߋ����� �����	��-�x�Q� c�u�������R�d�� B���	-?Q�� u�������� ��d��˰ew ����f��/ R+/=/O/a/s/�/, ��y�/�/�/�/?? )?�M?_?q?�/�?�? �?�?�?�?�/d�-��? ;OMO_OqO�O�O<?�O �O�O(O__%_7_I_ [_Od���O�_�_�_ �_�_o�O%o7oIo�_ moo�o�o�o�on_�W9So,>Pb 	os��Qo������(�:�ɪ	��0 �u���������Ϗv ����;�M�_�q� ����<�N�����9��  ��$�6�H��l�~� ��۟��Ưد���� ����ۥ�Z�l�~��� ����[�ؿ���G� � 2�D�V�h�z�!�[�n� ���������� �ǿ D�V�h߳όߞ߰��� ���ߍϟ���}�2�D� V�h�z��3߰����� ���
��.�@�R��� ��F����������� ����.@��dv ����e��Ų+U 
.@Rd� ������//<*/�  �	Y/ k/}/�/�/�/�/�/�/x�/?;   // 7/U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o�#<  
� (  ��M ( 	  �o�o�o�o�oC 1SUg����t��j?: �y *�<�N��r������� ��̏������a� >�P�b�t�����ߏ�� Ο��'���(�:�L� ^����������ʯܯ � ��$�k�}�Z�l� ~�ů����ƿؿ��� C� �2�Dϋ�h�zό� �ϰ���	�����
�Q� .�@�R�d�v߈����� ������)���*�<� N�`�߄������� ������&�m�J�\� n�������������� 3�E�"4F��j| ������ S0BTfx�� ����//,/ >/P/���/�/�/� �/�/�/??(?o/L? ^?p?�/�?�?�?�?�? �?5?O$O6O}?ZOlO�~O�O�O�O�?�p@ A�B�O�O_�C�G��`��#frh:�\tpgl\ro�bots\m10�iaAS_8l.xml�Oe_w_�_�_�_��_�_�_�_on�� o>oPoboto�o�o�o �o�o�o�oo: L^p����� �� ��6�H�Z� l�~�������Ə؏� ����2�D�V�h�z� ������ԟ���� 	�.�@�R�d�v����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶���������� XVA |�O+P<< )P ?���A���9�[� ��oߑ߿ߥ������� ���=�#�E�s�Y������������6��$TPGL_OUTPUT 1	A�	A !� -�B�T�f�x������� ��������,> Pbt�������-�!Є��2345678901 );M_g�2 ��������@/0/B/T/f/�}p/ �/�/�/�/�/x/�/? (?:?L?^?p??~?�? �?�?�?�?�?�?$O6O HOZOlOOO�O�O�O �O�O�O�O
_2_D_V_ h_z__�_�_�_�_�_ �_�_�_.o@oRodovo �o o�o�o�o�o�o �o<N`r� .������� "�J�\�n�����*����ȏڏ�������} �F�X�j�|��������@#�՟�)� ( 	 ��
�@� .�d�R���v������� �Я���*��N�<� ^���r�����̿��� ޿ ���J�8�n����8�vϨϺ͒��� �����$��
��U�g� �sߝ�w߉�����C� �����Q�c�=�� ���߁���i���� ��;�M���5�����/� ��������_�q�7 I��QYk�� %����3 i{���K�� ��///�/e/w/ /�/�/�/�/�/A/�/ ?+?�/O?a?;?M?�? �/?�?�?y?�?O�? OKO]O�?aO�O-OO �O�O�O�O_oO�OG_ �O3_}_�_i_�_�_#_ �_�_o�_1oCooOo yo�_�_�o�o[o�o�o �o�o-?�ocu�a�������)�WGL1.XM�L��(��$TPOFF_LIM ��|�����6��N_SV>�  ���P�P_MON7 2��R������22�STRT?CHK 3��P��C�9�VTCOM�PATe��T�VW�VAR 4��\�i� Ə *��I���:�_DE�FPROG %���%PART1 TLd�{���4��_DISPLAY�E���Z�INST_�MSK  �� ���INUSER�叜�LCK�QUICKMEN�ޜ�SCRE1������tpsc@���L�Q�P�b�_f��ST�P�RACE_CFG 5����I�	3�
?����HNL 26i�b�ѡ� ?��� )�;�M�_�q�������ITEM 27�� �%$1234567890ؿ�  =<���"�  !(�0�<��u�3�ֿ������ ��0���T�f�/ߊ�J� ��Z߀������4� >߸�b��4�F��j� ������l�������� ^������*�x��� �������6�H�l� ,��Pb��x��< � �D�(� 4���N��� �@ /dv�/$/ �~/�/��//*/�/ N/?r/2?D?�/Z?�/ �/�??�?&?�?�?~? n?�?�?�?�?0O�?�O �O�O"O�OFOXOjO�O �O:_`_r_�O~_�O_ _�_�_T_o&o�_2o �_�_�o�_�oo�o�o >o�obo�o=�oX�o h���(:L �p�B�T��x�� � �����6����l� �����k�Ə��ꏪ���� �ҟD�V����S�8��$��  ��$� ɡ{�r�
 ������үS��UD1:\߬���6�R_GRP �19Ż� 	 @{�*�<�&�\� J���n��������˿�ٺ��߯��'��?�  B�T�>�t�b� �φϼϪ�������� �:�(�^�L߂�pߒ߆��	�����4�S�CB 2:@� -�*�<�N�`�r������*�UTOR?IAL ;@�Ư��/�V_CONFIG <@�ġx��¯d��OUTPU�T =@�U���p�����������  2DVhz� R�������  2DVhz�� �����
//./ @/R/d/v/�/��/�/ �/�/�/??*?<?N? `?r?�?�?�/�?�?�? �?OO&O8OJO\OnO �O�O�?�O�O�O�O�O _"_4_F_X_j_|_�_ �O�_�_�_�_�_oo 0oBoTofoxo�o�o�_ �o�o�o�o,> Pbt���o�� ����(�:�L�^� p��������ʏ܏�  ��$�6�H�Z�l�~� ����>�P������� �(�:�L�^�p����� ������ܯ� ��$� 6�H�Z�l�~������� ůؿ���� �2�D� V�h�zόϞϰ���ӿ ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<�N�`�r�� ������������ &�8�J�\�n������� ����������"4 FXj|���� ����0BT fx������ �//,/>/P/b/t/ �/�/�/�/�/��/? ?(?:?L?^?p?�?�?�?�?�?������?�?�1�?&OɟJO \OnO�O�O�O�O�O�O �O�O_"_�/F_X_j_ |_�_�_�_�_�_�_�_ oo0oA_Tofoxo�o �o�o�o�o�o�o ,=oPbt��� ������(�9 L�^�p���������ʏ ܏� ��$�6�G�Z� l�~�������Ɵ؟� ��� �2�C�V�h�z� ������¯ԯ���
� �.�?�R�d�v����� ����п�����*� <�M�`�rτϖϨϺ� ��������&�8�I� \�n߀ߒߤ߶�����������"�4�C��$�TX_SCREE�N 1>�5;�0�}�C�� ��������u�2F t�!�3�E�W�i�{��� ������������� /��Sew��� $�H�+= O������� �V/z'/9/K/]/ o/�/��//�/�/�/ �/?#?�/�/Y?k?}? �?�?�?*?�?N?�?O�O1OCOUO�?yO�$�UALRM_MS�G ?c��p� qOFګO�O�O�O_ _6_)_;_Y___�_�_�_�_�_�ESEV � �M
f�BE�CFG @c��m�  F�@��  A:a   B�F�
 �_M�c� moo�o�o�o�o�o�o��o!/waGRPw 2A k 0F��	 Woy�@I_�BBL_NOTE� B jT���lM�h�O��,`�rDEFPRO��@%�K (%�PART2z�|% �_��?�*�c�N��� r��������̏��{�FKEYDATA� 1Cc�cpp 	/gF�fi�{�R�������,(���F�(POINT�z� ҐIREC��B�)�ND-�l�'�C?HOICE]p���TOUCHUP ����ȯ�ӯ���4� F�-�j�Q�������Ŀ�������ω����/frh/gu�i/whitehome.png)�`g�yϋϝϯπ@�pointR����ϰ��+ߺ�  A�direc��g�yߋ�8�߯�>�/inQ��������0��E�choicQ�o��������@�touchup_�����+��=���@�arwrg��w���������F� ���� $6H�� l~����U� � 2D�hz �����c�
/ /./@/R/�v/�/�/ �/�/�/_/�/??*? <?N?`?7�e?�?�?�? �?�?�?�/
OO.O@O ROdO�?�O�O�O�O�O �OqO�O_*_<_N_`_ r__�_�_�_�_�_�_ _o&o8oJo\ono�_ �o�o�o�o�o�o�o�o "4FXj|� �������0� B�T�f�x�������� ҏ������,�>�P� b�t��������Ο�� �����:�L�^�p�h����/����:���ۯ�8�ɯ�(��7�,�S��POINT\���Ϫ����ο��  CHOI�CE]��TOUCHUP��8� \�Cπ�gϤ϶ϝ��� �������4��X�j��Qߎ�m;��whitehom^��������������poinf�R�d�v��� %������������� <�N�`�r�������7�>5�choic�������'*�4�t?ouchup��e�w���,�4�arwrgA��� /2�Sew�� �<���//+/ =/�a/s/�/�/�/�/ J/�/�/??'?9?�/ ]?o?�?�?�?�?�?X? �?�?O#O5OGO�?kO }O�O�O�O�O��bO�O __1_C_U_\Oy_�_ �_�_�_�_b_�_	oo -o?oQoco�_�o�o�o �o�o�opo); M_�o����� ��~�%�7�I�[� m��������Ǐُ� z��!�3�E�W�i�{� 
�����ß՟����� �/�A�S�e�w���� ����ѯ������+� =�O�a�s���������Ϳ߿�Ϟ��}������:�@L�^�6πϒ�l�,~� ��v��������A� (�e�w�^ߛ߂߿��� �������+��O�6� s�Z��������� ��O'�9�K�]�o��� �������������� ��5GYk}� ������1 CUgy��,� ���	//�?/Q/ c/u/�/�/(/�/�/�/ �/??)?�/M?_?q? �?�?�?6?�?�?�?O O%O�?IO[OmOO�O �O�ODO�O�O�O_!_ 3_�OW_i_{_�_�_�_ @_�_�_�_oo/oAo �eowo�o�o�o�o�_ �o�o+=O�o s�����\� ��'�9�K��o��� ������ɏۏj���� #�5�G�Y��}����� ��şןf�����1� C�U�g����������� ӯ�t�	��-�?�Q� c�򯇿������Ͽ� 󿂿�)�;�M�_�q�  ϕϧϹ�������~� �%�7�I�[�m��V`����V`����߼��ݦ������,��3���W�>�{� ��t���������� ��/�A�(�e�L����� ����������  =$asRo��� ��� �'9K ]o����� ���#/5/G/Y/k/ }//�/�/�/�/�/�/ ?�/1?C?U?g?y?�? ?�?�?�?�?�?	O�? -O?OQOcOuO�O�O(O �O�O�O�O__�O;_ M___q_�_�_$_�_�_ �_�_oo%o�_Io[o moo�o�o2o�o�o�o �o!�oEWi{ �������� �/�6S�e�w����� ����N������+� =�̏a�s��������� J�ߟ���'�9�K� ڟo���������ɯX� ����#�5�G�֯k� }�������ſ׿f��� ��1�C�U��yϋ� �ϯ�����b���	�� -�?�Q�c��χߙ߫� ������p���)�;� M�_��߃������h�����p����p����,�>��`�r�L�,^��V ����������!E W>{b���� ���/S: w�p����� //+/=/O/a/p�/ �/�/�/�/�/�/�/? '?9?K?]?o?�/�?�? �?�?�?�?|?O#O5O GOYOkO}OO�O�O�O �O�O�O�O_1_C_U_ g_y__�_�_�_�_�_ �_	o�_-o?oQocouo �oo�o�o�o�o�o �o);M_q�� $������� 7�I�[�m���� ��� Ǐُ����!��E� W�i�{�������ß՟ �����/���S�e� w�������<�ѯ��� ��+���O�a�s��� ������J�߿��� '�9�ȿ]�oρϓϥ� ��F��������#�5� G���k�}ߏߡ߳��� T�������1�C��� g�y��������b� ��	��-�?�Q���u� ����������^���@);M_6�a��6������������, ��7[mT �x�����/ !//E/,/i/{/b/�/ �/�/�/�/�/�/?? A?S?2�w?�?�?�?�? �?���?OO+O=OOO aO�?�O�O�O�O�O�O nO__'_9_K_]_�O �_�_�_�_�_�_�_|_ o#o5oGoYoko�_�o �o�o�o�o�oxo 1CUgy�� ������-�?� Q�c�u��������Ϗ �����)�;�M�_� q��������˟ݟ� ���%�7�I�[�m�� ��h?��ǯٯ���� �3�E�W�i�{����� .�ÿտ����Ϭ� A�S�e�wωϛ�*Ͽ� ��������+ߺ�O� a�s߅ߗߩ�8����� ����'��K�]�o� �����F������� �#�5���Y�k�}��� ����B������� 1C��gy��� �P��	-? �cu�����ڦ���������/-�@/R/,&,>?�/6?�/�/ �/�/�/?�/%?7?? [?B??�?x?�?�?�? �?�?O�?3OOWOiO PO�OtO�O�O���O�O __/_A_Pe_w_�_ �_�_�_�_`_�_oo +o=oOo�_so�o�o�o �o�o\o�o'9 K]�o����� �j��#�5�G�Y� �}�������ŏ׏� x���1�C�U�g��� ��������ӟ�t�	� �-�?�Q�c�u���� ����ϯ�󯂯�)� ;�M�_�q� ������� ˿ݿ���O%�7�I� [�m�φ��ϵ����� ����ߞ�3�E�W�i� {ߍ�߱��������� ��/�A�S�e�w�� ��*���������� ��=�O�a�s�����&� ��������'�� K]o���4� ���#�GY k}���B�� �//1/�U/g/y/ �/�/�/>/�/�/�/	?�?-???�A;�>����j?|? �=f?�?�?�6,�O�? �OO�?;OMO4OqOXO �O�O�O�O�O�O_�O %__I_[_B__f_�_ �_�_�_�_�_�_!o3o �Woio{o�o�o�o�/ �o�o�o/A�o ew����N� ���+�=��a�s� ��������͏\��� �'�9�K�ڏo����� ����ɟX�����#� 5�G�Y��}������� ůׯf�����1�C� U��y���������ӿ �t�	��-�?�Q�c� �ϙϫϽ�����p� ��)�;�M�_�q�Ho �ߧ߹���������� %�7�I�[�m���� �����������!�3� E�W�i�{�
������� ��������/AS ew����� ��+=Oas ��&����/ /�9/K/]/o/�/�/ "/�/�/�/�/�/?#? �/G?Y?k?}?�?�?0? �?�?�?�?OO�?CO�UOgOyO�O�O�O����K�������O�O�M�O _2_V,oc_o�_n_�_�_ �_�_�_oo�_;o"o _oqoXo�o|o�o�o�o �o�o�o7I0m T�������� �!�0OE�W�i�{��� ����@�Տ����� /���S�e�w������� <�џ�����+�=� ̟a�s���������J� ߯���'�9�ȯ]� o���������ɿX�� ���#�5�G�ֿk�}� �ϡϳ���T������ �1�C�U���yߋߝ� ������b���	��-� ?�Q���u����� ������)�;�M� _�f������������ ��~�%7I[m ��������z !3EWi{
 �������/ //A/S/e/w//�/�/ �/�/�/�/?�/+?=? O?a?s?�??�?�?�? �?�?O�?'O9OKO]O oO�O�O"O�O�O�O�O �O_�O5_G_Y_k_}_ �__�_�_�_�_�_o�o�$UI_IN�USER  ����@a��   o$o_�MENHIST �1D@e � ( M`���(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153�,1_o�o�o�o�9)�o�o422�oU�gy�,xedi=t�bMAIND�8��� �'�/~71�[�m�����Q�o6�154J�������P��>�P�b� t�����'���Ο��� ����:�L�^�p��������4��a4�ѯ� ����+�.�O�a�s� ������8�Ϳ߿�� �'϶�ȿ]�oρϓ� �Ϸ�F��������#� 5���Y�k�}ߏߡ߳� B�T�������1�C� ��g�y�����אָ ����	��-�?�Q�T� u�����������^��� );M_��� �����l %7I[��� ����z/!/3/ E/W/i/��/�/�/�/ �/�/����?/?A?S? e?w?z/�?�?�?�?�? �?�?O+O=OOOaOsO �OO�O�O�O�O�O_ �O'_9_K_]_o_�__ �_�_�_�_�_�_o�_ 5oGoYoko}o�oo�o �o�o�o�o�/
?C Ugy���o�� ��	����Q�c� u�������:�Ϗ�� ��)���M�_�q��� ����6�H�ݟ��� %�7�Ɵ[�m������ ��D�ٯ����!�3����$UI_P�ANEDATA �1F���i��  	��}  frh/c�gtp/flex�dev.stm?�_width=0�&_height�=10����ice�=TP&_lin�es=15&_c�olumns=4���font=24�&_page=w�hole��E�!v)�  rim��  z�(�:�L�^�pς� 鿔ϸϟ����� �� ��6��Z�l�Sߐ�w����߭���!v� ��     ��"�}���J��2��39ཾ1ϵ/doub*�2���ual���$����� ����/���S�:�w� ��p����������� ��+OaH����
�   �i������ %xI��m� ���.���!/ /E/W/>/{/b/�/�/ �/�/�/�/�/?/?�I6k�fk?}?�?�? �?�??�?\OO1O COUOgO�?�O�O�O�O �O�O�O�O__?_&_ c_u_\_�_�_�_�_B? T?oo)o;oMo_o�_ �o�?�o�o�o�o�o zo7[B� x������� 3�E�,�i��_�_���� ÏՏ���L��/��o S�e�w��������џ ������+��O�a� H���l�������߯Ư �v���F�K�]�o��� ������ɿ<����� #�5�GϮ�k�}�dϡ� �����Ͼ������� C�U�<�y�`ߝ߯�"� 4�����	��-�?�� c�ֿ��������� ��Z����;�"�_�q� X���|�����������@%I�����T@������){ ��8J\n� �������/ �4//X/j/Q/�/u/��/�/�/�/x�������$UI_POST�YPE  ���� 	 ��/K?2QUICK�MEN  );�8?N?0RESTO�RE 1G���  ��*defaul�tx�DOUB�LE�=DUA�L�?medit�page,PART1,1�?*O<ONO|`OBmenuB154O�O�O�O�O �6�O�O__/_A_�1 �/R_d_�O�_�_�_�_ �_�_�_o/oAoSoeo o�o�o�o�o�o|_�o �oto=Oas� (������� '�9�K�]�o�|��� ���ۏ����#�Ə G�Y�k�}���2���ş ן��������,��� P�y���������d�� ��	��-�ЯQ�c�u�x����S=SCREi0�?n=u1�sc�0u2ڴ3�ڴ4ڴ5ڴ6ڴ7rڴ8ڱ��TAT%=�� }3��:UScER����Ӵksܳ�m�3m�4m�5m�6�m�7m�8m�0ND�O_CFG H�);d c0PD��W��Non�e\2N�_INFOW 1I���{00%���x�
�K�.� o߁�dߥ߷ߚ��߾� �����5�G�*�k�R<���OFFSET L)9�x�@��0 H�����������(� U�L�^���b������� ������$6��~?�p�
����_UFRAM�0@������RTOL_�ABRT���E�NB GRP �1M�9z1Cz  A�ec��cu ������h0�U/��MSK � 2�N��%���%Rs/ _'EVN2$�ƈ&v��2N��
 h���UEV!�td:\event_user\w/F� C7�/�B�F<��!SP�!�'sp�otweld=!C6????�0b$!b/�/�?�?�7!�? �?�?OAO�?�?wO"O �OFOXOjO�O�O_�O �O�OO_>_s__0_f_ �_�_�_�_�_o�_9o Ko�_o�o,o�oPobj~�&WRK 2OX�F�8�o	 �o @R-v�c�� �����*��N� `�;�����q���̏���ݏ���$VARS_CONFI���P�� FP@����CCRG��SP��Z@�9�D��B�BH�p����Ce���їϑ?�ᐶU�MRK2Y��)B�	��C�X��1: SC13?0EF2 *3�7��@����ch �5�B����A@��C�Ȑ� ��� ��9���ȯ�����"���ӑ��	�Z���� B��� u���z����᯾��� �Ϳ��*��'�`� ��Aϖρϓ������\�X�TCCc�ZR��4��pa��'�G�F,��![�� ��a 2345678901q�y�'9�n���n߰ߘ#����j�$����B��Ӗ ��ϑ?:�o=L{�� !p� �p��ia/[�� �Ԇ���������� )�;�(�:�q��p��� ���������%� I�[�H���{���������"�S�SELE�C�$!?�AVIoA_WO�`\T)�_ff,		��= �;G�P ��R'	�RTSYN'CSE�j��n�e�WINURL ?u��R����� //"�ISI�ONTMOU�/ ��*%c�]S۳��S۵@/� �FR:\,#\D�ATAs?MЄ� wMCk&LOGx/   UD1k&�EX�/��' ?B@ ���"�!�DESKTOP�-MC6FJ6K��/�#?%?�le �� n6  �����f�"�� -��N5K�   =���w1��t0� }�(TRAIN�/hH҆2�bd�3pw5>{4 #`�"'(:��^]� (���9 M��OO+O=OOO�O sO�O�O�O�O�O�O�O�_$(STAT _'� �z�b_t_�_�hq$�_�_'%_GES#�`]���0 �
����R�WHOMI}NV aS۾�`��b"���C�ז�&�WJMPERR� 2b]�
   =�jho^l��o�o�o �o�o�o�o.<�m`r�S_� R�EV cO^#�LEXr�Td7��1-e�_�VMPHASE � j���&�O�FFo_ENB � \�	P2R$e/SۿN��c|3�@:�`Q�u����?s33�4�1K� g�']g�t�g��&�S`�hWm�3�\BQ���C�F����81��_�
�A/�4��/�7k� B��C.�\@�4��� S�4�0�3��o�=�,������5ǟ[�s�C�;��Ԙ�#��rͫSAq��9��;�M�����Cj��ԓ�l��+&eB\�%�ՀS���_�u���������]�o��+��������%���6��+F�h_�����A�W������^Cr �B��+T�������*�dC�	Ml߯Կ�M�C�LA;B�6x��i敚,2��3��*ȹO��a�7�1�{�p������cda*�9�ӯɿ���C �����x�m�'�Y�K�	��e�Z����A�AC����Փ#�Ln��2A����Ϝ�����:6�B�������+�B)m�)�����C߀8�X��߄�� [��������3� ���i�^�p������ ������� /�!S� Hw�����y��� ���+=2a��_q��ÅTD�_FILTES`i��[ Է��P�� <//'/9/K/]/o/ �/�/�/6��/�/�/ ??,?>?P?b?t?�Y�SHIFTMENoU 1jWm<�|%��?�t�?�?O�? �?EOO.O{OROdO�O �O�O�O�O�O�O/__�	LIVE/S�NAP#Svsf�liv�~A_�^�PION &�U^PdRmenuz___��_�_�r�5G�kΉ�ֈ9MOG�l�~�z�łZDdm��a<�ۀ �P�$WA�ITDINEND�  �U��#bxfO9K-��oOUT�o�h�S�o�iTIM�e���lGo}�o2{��oz�oz�o�hREcLE�.��hTM^{�d�xc_ACT�WP-���h_DATA n΅�N�3�<E��RDIS�P�~��$XVRa�o9n�$ZABC_GRP 1p[k ,2J��=Qa��pVSPT q�9m���
�Z��_��Z)�?�އDCSCH`r#�����[IPbs[o!�۟���؊MPCF__G 1t����A0� O����u���Ġp�� 	�?���o`�  ?���2?�k��1�?�ɾ�����4/6��u��D5Oy���C���?����<� ���>%��6�����u=C������ί�1� ���	������˿� � 8��h�Ca���.~:��1�G�����۸��� &� �2�H�Vπ��,�>��0V�h��� �`�v����_CYLI�ND�w(� ��� ,(  * E�V��B��fߣߊ� ��������?� � ��D�+�=�z�ߞ�� ������g���@��'���v����̞�2x �� �=���? ��	��-=��`��zA��SPH�ERE 2y%�� ��*����X� kFX��|� ���///ew T/�x/_/q/�/��/��/�/��ZZ�v � f