��  I��A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����SBR_T �  | 	$S�VMTR_ID � $ROBO�T9$GRP�_NUM<AXIaSQ6K 6NFF�3 _PARAM�F	$�  �,$MD SPD�_LIT��&2�*  � ��  ��$$C�LASS  ����������� VERSION��  ���IRTUAqL��'  1 �� T����ARC Mat�e 100iC/�8���  �aiS8/400�0 40A��
�H1 DSP1-�S1��	P01�.03W,  �	�  ��PCR �� �C������0��
=��0�r9  �3!M�����  H� � �"`��� ���  k ���~Z yy������C�W�� 1�3����?$�p��B:o~�L����&�����P ���7� H���������g u � y���e���%��.���fB�� � d� ��c ��8 :?����'b:
�c/�/�/�/?��3?;?f<?a?�s?�?��1�1���>�������q��2��%��0*�G��"�DJ���?�?"4p<N`r2|2�����@��{vA�@?}9}��� ������X � %p��1#� ��� 3�|��=�'���r� ���:+����� ��'�� sBZ ��?��d%z'	?��8U�'��/�/�D �/�_�_�_�_!?�_E?�o o2oDo 1�2����?�� �\p �	< ��2.���>���� d� ��	� ��o�o�m�?NB2/5
 A2m3|GB@ORE;
� �  V@�������wD� ��<��9"�b8 lѿ  ���E&���4�&"m"īa" �0~#�0�3�B\`�( ��] �qC��:+�� ��/�� TV$��o�� �  2|!���-�"�pHX�c9	`�� # (���� ��jTqrYa�J�\�n����_ ���_ȏڏ����"��4�F���P�oN�biS0.5S/6�kx4|4�o�NIp�ϓ ��7_�K����2���p�����DsFp 8z ��������o�	��]!�$��S@A�S���o.�r� +V$�b��o9 ]�s;T@�;�����}�T��2pr���"��rY�ZP���
	���#�5� ��Y���}�������ſ׿�����Rh�R���R��x5�|5����О�����<<l���@�
b��� ,�>���? �����rZ 1�@�n���9�s�X@g��x�e�DJV ïկ���������A� 
�e�w�@�R�d�v��8���� ��NU@�4I�6|6d��{@��d�R�a���8tG�8��a�Sn�Ҵ��
�8��]����Ͻ����� �N �� �2Z �����tX���s�  ��1���D|ߎؐrY �}���� t��� ��� ��$����#5GYk�
�?����x��(���7�	�t����/ /2/D/ V/h/z/�/�/�/�/�/��/�/
??.?@?P<� P?t?�?�?�?�?�?�? �?OO(O0C��FO ����O�O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_o^? &o8oJo\ono�o�o�o �o�o�o6OhOZO#~O �OXj|���� �����0�B�T� f�x�������
o��� ����,�>�P�b�t� �����o����*<N �(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�ȏ������ ƿؿ���� �2�D� V�ҟğn������� ����
��.�@�R�d� v߈ߚ߬߾������� ��*N�`�r�� �����������^� �ς�K��ϸπ����� ����������"4 FXj|���� �2��0BT fx������ �R�d�v�>/P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? ��?�?�?�? OO$O 6OHOZOlO~O���O /"/4/�O_ _2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRo�? vo�o�o�o�o�o�o�o *�O�O�Os�O �O������� &�8�J�\�n������� ��ȏڏ���Zo�4� F�X�j�|�������ğ ֟�D� �z�� f�x���������ү� ����,�>�P�b�t� ������������ �(�:�L�^�pςϔ� ��"����8�J�\�$� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z�ֿ������� ����
��.�@�R��� ���ϛ���������� *<N`r� ������ &��8\n��� �����/l�5/ (/�������/�/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? @OO,O>OPObOtO �O�O�O�O�OJ/</�O `/r/�/L_^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�? �o�o�o�o 2D Vhz�O_�O�_ 0_�
��.�@�R�d� v���������Џ�� ��*�<�N��o`��� ������̟ޟ��� &�8��]�P���� ��ȯگ����"�4� F�X�j�|�������Ŀ ֿ����h�0�B�T� f�xϊϜϮ������� ��r�d�߈�����t� �ߘߪ߼�������� �(�:�L�^�p��� �����&��� ��$� 6�H�Z�l�~������� 0�"���F�X� 2D Vhz����� ��
.@Rd v������� //*/</N/`/���/ x/���/�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O �XOjO|O�O�O�O�O �O�O�O__�/�/6_ �/�/�/�_�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�oNO (:L^p�� ���&_X_J_�n_ �_H�Z�l�~������� Ə؏���� �2�D� V�h�z������o��ԟ ���
��.�@�R�d� v���������,�>� ��*�<�N�`�r��� ������̿޿��� &�8�J�\ϸ��ϒϤ� �����������"�4� F�¯��^�د����� ��������0�B�T� f�x���������� ����v�>�P�b�t� ��������������N� ��r�;�ߨ�p�� ����� $ 6HZl~��� �"���/ /2/D/ V/h/z/�/�/�/�/ �/BTf.?@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O ��O�O�O�O�O__ &_8_J_\_n_�/�/�_  ??$?�_�_o"o4o FoXojo|o�o�o�o�o �o�o�o0B�O fx������ ���v_�_�_c��_ �_������Ώ���� �(�:�L�^�p����� ����ʟܟ�J �$� 6�H�Z�l�~������� Ưد4����j�|��� V�h�z�������¿Կ ���
��.�@�R�d� vψϚϬ�������� ��*�<�N�`�r߄� ������(�:�L�� &�8�J�\�n���� �����������"�4� F�X�j��ώ������� ������0B�� ���ߋ������� �,>Pbt �������/ /r�(/L/^/p/�/�/ �/�/�/�/�/ ?\%? ?���~?�?�?�? �?�?�?�?O O2ODO VOhOzO�O�O�O�O�O 0/�O
__._@_R_d_ v_�_�_�_�_:?,?�_ P?b?t?<oNo`oro�o �o�o�o�o�o�o &8J\n���O ������"�4� F�X�j��_�_�_��o  o�����0�B�T� f�x���������ҟ� ����,�>��P�t� ��������ί��� �(���M�@���̏ޏ ����ʿܿ� ��$� 6�H�Z�l�~ϐϢϴ� ��������X� �2�D� V�h�zߌߞ߰����� ��b�T���x�����d� v����������� ��*�<�N�`�r��� ����������� &8J\n����  ���6�H�"4 FXj|���� ���//0/B/T/ f/��x/�/�/�/�/�/ �/??,?>?P?�u? h?���?�?�?O O(O:OLO^OpO�O�O �O�O�O�O�O __$_ �/H_Z_l_~_�_�_�_ �_�_�_�_o�?|?&o �?�?�?�o�o�o�o�o �o�o
.@Rd v������>_ ��*�<�N�`�r��� ������oHo:o�^o po8�J�\�n������� ��ȟڟ����"�4� F�X�j�|������į ֯�����0�B�T� f�x�ԏ����
��.� ����,�>�P�b�t� �ϘϪϼ�������� �(�:�Lߨ�p߂ߔ� �߸������� ��$� 6ﲿ��N�ȿڿ쿴� ��������� �2�D� V�h�z����������� ����
f�.@Rd v������>� p�b�+���`r� ������// &/8/J/\/n/�/�/�/ �/�/�/�/?"?4? F?X?j?|?�?�?��? �?2DVO0OBOTO fOxO�O�O�O�O�O�O �O__,_>_P_b_t_ �/�_�_�_�_�_�_o o(o:oLo^o�?�?vo �?OO�o�o $ 6HZl~��� ����� �2��_ V�h�z�������ԏ ���
�fo�o�oS��o �o��������П��� ��*�<�N�`�r��� ������̯ޯ:��� &�8�J�\�n������� ��ȿ$���Z�l�~� F�X�j�|ώϠϲ��� ��������0�B�T� f�xߊߜ��������� ����,�>�P�b�t� ��������*�<�� �(�:�L�^�p����� ���������� $ 6HZ��~��� ���� 2�� ���{������ ��
//./@/R/d/ v/�/�/�/�/�/�/�/ ?b?<?N?`?r?�? �?�?�?�?�?�?LO O���nO�O�O�O �O�O�O�O�O_"_4_ F_X_j_|_�_�_�_�_  ?�_�_oo0oBoTo foxo�o�o�o*OO�o @OROdO,>Pbt �������� �(�:�L�^�p����_ ����ʏ܏� ��$� 6�H�Z��o�o�o���o ؟���� �2�D� V�h�z�������¯ԯ ���
��.���@�d� v���������п��� ��t�=�0Ϫ���Ο �ϨϺ��������� &�8�J�\�n߀ߒߤ� ��������H��"�4� F�X�j�|������ ��R�D���h�zό�T� f�x������������� ��,>Pbt ������� (:L^p��� ���&�8� //$/ 6/H/Z/l/~/�/�/�/ �/�/�/�/? ?2?D? V?�h?�?�?�?�?�? �?�?
OO.O@O�eO XO����O�O�O�O __*_<_N_`_r_�_ �_�_�_�_�_�_oo p?8oJo\ono�o�o�o �o�o�o�o�ozOlO �O�O�O|���� �����0�B�T� f�x���������ҏ.o ����,�>�P�b�t� ������8*�N `(�:�L�^�p����� ����ʯܯ� ��$� 6�H�Z�l�~�ڏ���� ƿؿ���� �2�D� V�h�ğ�π����� ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<`�r�� ������������ &��ϔ�>������Ϥ� ����������"4 FXj|���� ���V�0BT fx�����.� `�R�/v���P/b/t/ �/�/�/�/�/�/�/? ?(?:?L?^?p?�?�? �?�?�?�? OO$O 6OHOZOlO~O�O��O �O"/4/F/_ _2_D_ V_h_z_�_�_�_�_�_ �_�_
oo.o@oRodo �?�o�o�o�o�o�o�o *<N�O�Of �O�O_����� &�8�J�\�n������� ��ȏڏ����"�~o F�X�j�|�������ğ ֟���V�zC�� �x���������ү� ����,�>�P�b�t� ��������ο*��� �(�:�L�^�pςϔ� �ϸ������J�\�n� 6�H�Z�l�~ߐߢߴ� ��������� �2�D� V�h�z��述����� ����
��.�@�R�d� v����ώ���,��� *<N`r� ������ &8J��n��� �����/"/~� ����k/�����/�/�/ �/�/�/??0?B?T? f?x?�?�?�?�?�?�? �?RO,O>OPObOtO �O�O�O�O�O�O</_ �Or/�/�/^_p_�_�_ �_�_�_�_�_ oo$o 6oHoZolo~o�o�o�o O�o�o�o 2D Vhz��__� 0_B_T_�.�@�R�d� v���������Џ�� ��*�<�N�`�r��o ������̟ޟ��� &�8�J�������  �ȯگ����"�4� F�X�j�|�������Ŀ ֿ�����z�0�T� f�xϊϜϮ������� ���d�-� ߚ����� �ߘߪ߼�������� �(�:�L�^�p��� �������8� ��$� 6�H�Z�l�~������� ��B�4���X�j�|�D Vhz����� ��
.@Rd v������� //*/</N/`/r/��  ���/(�/?? &?8?J?\?n?�?�?�? �?�?�?�?�?O"O4O FO�XO|O�O�O�O�O �O�O�O__0_�/U_ H_�/�/�/�_�_�_�_ �_oo,o>oPoboto �o�o�o�o�o�o�o `O(:L^p�� �����j_\_� �_�_�_l�~������� Ə؏���� �2�D� V�h�z������� ���
��.�@�R�d� v������(���>� P��*�<�N�`�r��� ������̿޿��� &�8�J�\�n�ʟ�Ϥ� �����������"�4� F�Xߴ�}�p����� ��������0�B�T� f�x���������� ����,���P�b�t� �������������� �߄�.�ߺ��ߔ ����� $ 6HZl~��� ���F�/ /2/D/ V/h/z/�/�/�/�/ PB?fx@?R?d? v?�?�?�?�?�?�?�? OO*O<ONO`OrO�O �O��O�O�O�O__�&_8_J_\_n_�_�%��$SBR2 1� 5�P T0? �  C?7 �_�_�_o o2oDo Vohozo�o�o�o�o�o�Q�o�_!3E Wi{����� ���o� A�S�e� w���������я�����+��5�.�o� ��������ɟ۟��� �#�5�G�Y�<�}�`� ����ůׯ����� 1�C�U�g�y���n��� ��ӿ���	��-�?� Q�c�uχϙϫϽ��~�_�����!�3�E� W�i�{ߍߟ߱����� �������(�:�L�^� p�����������  �����H�Z�l�~� ��������������  2D(�:�z�� �����
. @RdvZ��� ���//*/</N/ `/r/�/�/�/��/�/ �/??&?8?J?\?n? �?�?�?�?�?�?�/�? O"O4OFOXOjO|O�O �O�O�O�O�O�O_�? 0_B_T_f_x_�_�_�_ �_�_�_�_oo,o>o "_boto�o�o�o�o�o �o�o(:L^ pTo������  ��$�6�H�Z�l�~� �����Ə؏����  �2�D�V�h�z����� ��������
��.� @�R�d�v��������� Я���؟�*�<�N� `�r���������̿޿ ���&�
�4�\�n� �ϒϤ϶��������� �"�4�F�X�<�|ߎ� �߲����������� 0�B�T�f�x��n߮� ����������,�>� P�b�t����������� ����(:L^ p������� ��$6HZl~ �������/  /D/V/h/z/�/�/ �/�/�/�/�/
??.? @?R?6/v?�?�?�?�? �?�?�?OO*O<ONO `OrOV?h?�O�O�O�O �O__&_8_J_\_n_ �_�_�_�O�O�_�_�_ o"o4oFoXojo|o�o �o�o�o�o�_�o 0BTfx��� ������o,�>� P�b�t���������Ώ �����(�:��^� p���������ʟܟ�  ��$�6�H�Z�l�P� ������Ưد����  �2�D�V�h�z����� ��¿Կ���
��.� @�R�d�vψϚϬϾ� �ϴ�����*�<�N� `�r߄ߖߨߺ����� �����&�8�J�\�n� ������������� �"���X�j�|��� ������������ 0BT8�J���� ����,> Pbt�j��� ��//(/:/L/^/ p/�/�/�/�/��/�/  ??$?6?H?Z?l?~? �?�?�?�?�?�?�/O  O2ODOVOhOzO�O�O �O�O�O�O�O
__ O @_R_d_v_�_�_�_�_ �_�_�_oo*o<oNo 2_ro�o�o�o�o�o�o �o&8J\n �do������ �"�4�F�X�j�|��� �����֏����� 0�B�T�f�x������� ��ҟ��ȏ��,�>� P�b�t���������ί ������:�L�^� p���������ʿܿ�  ��$�6��D�l�~� �Ϣϴ����������  �2�D�V�h�Lόߞ� ����������
��.� @�R�d�v���~߾� ��������*�<�N� `�r������������� ��&8J\n �������� ��"4FXj|� ������// 0/T/f/x/�/�/�/ �/�/�/�/??,?>? P?b?F/�?�?�?�?�? �?�?OO(O:OLO^O pO�Of?x?�O�O�O�O  __$_6_H_Z_l_~_ �_�_�_�O�O�_�_o  o2oDoVohozo�o�o �o�o�o�o�_�o. @Rdv���� ������o<�N� `�r���������̏ޏ ����&�8�J�.�n� ��������ȟڟ��� �"�4�F�X�j�|�`� ����į֯����� 0�B�T�f�x������� ��ҿ�����,�>� P�b�tφϘϪϼ��� ��Ŀ��(�:�L�^� p߂ߔߦ߸�������  ����6�H�Z�l�~� �������������  �2��(�h�z����� ����������
. @RdH�Z���� ���*<N `r��z��� �//&/8/J/\/n/ �/�/�/�/�/��/�/ ?"?4?F?X?j?|?�? �?�?�?�?�?�?�/O 0OBOTOfOxO�O�O�O �O�O�O�O__,_O P_b_t_�_�_�_�_�_ �_�_oo(o:oLo^o B_�o�o�o�o�o�o�o  $6HZl~ �to������  �2�D�V�h�z����� ������
��.� @�R�d�v��������� П�Ə؏�*�<�N� `�r���������̯ޯ �����
�J�\�n� ��������ȿڿ��� �"�4�F�*�T�|ώ� �ϲ����������� 0�B�T�f�x�\Ϝ߮� ����������,�>� P�b�t������� ������(�:�L�^� p���������������  $6HZl~ ������� ��2DVhz�� �����
//./ @/$d/v/�/�/�/�/ �/�/�/??*?<?N? `?r?V/�?�?�?�?�? �?OO&O8OJO\OnO �O�Ov?�?�O�O�O�O _"_4_F_X_j_|_�_ �_�_�_�O�O�_oo 0oBoTofoxo�o�o�o �o�o�o�o�_,> Pbt����� ����(�L�^� p���������ʏ܏�  ��$�6�H�Z�l�