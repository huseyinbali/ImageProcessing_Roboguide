��   v��A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@��?&�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	��&USRVI| 1  < `��R*�R��QPRIƍm� t1�PTR�IP�"m�$$C�LASP ��)�a��R��R `\ �SI�	g�  �aIR�Ts1	o`'2 L1���L1���R	 �,��?����a1`�b�ba� ����y`��  ����
 ��a�o�o1CU �oz�� ���c�
��.� @�R��v��������� Џ�q���*�<�N� `��������̟ޟ m���&�8�J�\�n� ��������ȯگ�{� �"�4�F�X�j����������Ŀֿ���`�TPTX��p���/�` s����$/soft�part/gen�link?hel�p=/md/tpmenu.dg�� �ϨϺ��υ����� &�8�J���n߀ߒߤ� ����W������"�4� F�X���|�����������a�f8�b�b�� ($p�-�@���T�?�x���a��a��c���c���� l���c��ah�a�h�h�2�h�	.f��������q�`���`  ���|f ep��*h#h�Fd��g�Xc�B 1)hR �\ _� �REG VE�D]���who�lemod.ht}m�	singl	�doub �trip8browsQ��� ��u���//�@/���dev�.sl�/3� 1�,	t�/_�/;/i/ ??/?�/S?e?w?�?�?�?� H`�?�?  OO$O6OHOZOlO~O�F @�?�O�O�O�O �O_�F�	�?�?;_M_ __q_�_�_�_�_�_�_ �_oo%o7oIo[omo oM'�o�o�o�o�o�o +=Oas� ��������? >�P�b�t��������� Ώ���O�����L� ^�_'_�������ş �����6�1�C�U� ~�y�����Ư��ӯ�o ���-�?�Q�c�u� ��������Ͽ��� �)�;�M�_�-��Ϭ� ����������*�<� 7�`�r�A�Sߨߺ�q� ��i�����!�J�E� W�i��������� ����"��/���O�I� w��������������� +=Oas� ������, >Pbt���߼ ���//����� ^/Y/k/}/�/�/�/�/ �/�/�/?6?1?C?U? ~?y?�?Y��?�?�?�? �?	OO-O?OQOcOuO �O�O�O�O�O�O�O_ _�R_d_v_�_�_�_ �_�_�_�_�o*o�_�o`oro�j�$UI�_TOPMENU� 1K`�aR 
d�a�*Q)*defa�ult5_]*�level0 * [	 �o�0��o'rtpio�[23]�8tpst[1[x)w9��o	�=h58E�01_l.png���6menu5�y�p�13�z��zb	�4���q��]� ��������̏ޏ)Rr����+�=�O�a����prim=�pa�ge,1422,1h�����şן����1�C�U�g����|�class,5�p�����ɯۯ�����13��*�<�N�`�4r���|�53�������ҿ�����|�8 ��1�C�U�g�y�����@����������"Y�` �a�o/��m!ηq�Y���avtyl}Tfqm�f[0nl�	��c�[164[w��59`[x�qG�y��tC8�|�29��o�%�1�� �{��m��!����� 0�B���f�x���������o���80�� '9K~���2P� ����\�� '9K����� �������1��/�$/6/H/Z/U�|�ainedi'ߑ/�/�/�/�/P�con�fig=sing�le&|�wintp���/$?6?H?Z?!Z �a�h?�?�e�?�� �?�?�?OO+O=OOO �?[O�O�O�O�O�O�O �O_a�%_L_^_p_�_ �_�_U��_�_�_ oo $o�_HoZolo~o�o�o 1o�o�o�o�o 2 �oVhz���? ���
��.��@� d�v���������M�� ���*�<�ˏ`�r� ��������^��;�M�sc���;���s �� �}���e�u��X��@�F7L���`��t꒯4�j�X�6e�u7�����ｿϿ������27��G�Y� k�}Ϗ��0�s����P�����!�1� M�_�q߃ߕ�T����� �������7�I�[� m����������� ���!�����6(�]��o��������$��74 6�����)t<ϯ�\�5	TPTX[�209©|Dw24`§J��
�w18�@�� ����0�2��A#��[	�t�v`�RxL�u1E0�1���5S:�$�treeview�3��3��&dua�l=o'81,26,4�O/a/s/2� �/�/�/�/�/�/�/?@'?9?K?]?o?��;/&�3$/6$���?�?�? 
?#O5OGOYOkO}O�?$�? "2�?8"2K��O�O_�O��1�?�E�Ϙg_y_�_�6_��edit��>_P_�_�_ o��/���_�Cooo �o�oB�o�o��oA �o�+=Oa s��o����� ��(�9���Q�x��� ������ҏO���� ,�>�P�ߏt������� ��Ο]�����(�:� L�^�ퟂ�������ʯ ܯk� ��$�6�H�Z� �l�������ƿؿ� y�� �2�D�V�h��� �Ϟϰ������ϕo�o ��o@ߧE�c�u߇� �߽߬�����O���� )�<�M�_�q���W� ��������&�8��� \�n���������E��� ����"4��Xj |����S�� 0B�fx� ���O��// ,/>/P/�t/�/�/�/ �/�/]/�/??(?:? L?��߂?1ߦ?�� �?�?�?�?O$O5OGO �?SO}O�O�O�O�O�O �O�O��2_D_V_h_z_ �_�_�/�_�_�_�_
o o�_@oRodovo�o�o )o�o�o�o�o* �oN`r���7 �����&��J� \�n���������E�ڏ ����"�4�ÏX�j� |�������a?s?蟗? �sO_/�A�S�e�w� ������������� �,�=�O�a�#_���� ��ο��=��(�:� L�^�pς�Ϧϸ��� ���� ߏ�$�6�H�Z� l�~�ߐߴ������� ����2�D�V�h�z� ������������
� ���@�R�d�v����� )���������ƚ�Ԕ*defau�lt%��*level8�ٯw����? tpsOt[1]�	�y��tpio[23���u���J�\menu7__l.png_|13��5�{�y4�u6���/ /'/9/K/]/���/�/ �/�/�/�/j/�/?#?�5?G?Y?k?�"pr�im=|page,74,1p?�?�?��?�?�?�"�6cl?ass,13�?*O@<ONO`OrOOB5xO@�O�O�O�O�O�#L �O0_B_T_f_x_{?�218�?�_�_�_�_�__B6o9oKo]ooo��o`�$UI_U�SERVIEW �1֑֑R 
���o��o�o[m�o' 9K] ���� �l���#�5��o B�T�f������ŏ׏ 鏌���1�C�U�g� 
���������ӟ~��� ��v�?�Q�c�u��� *�����ϯ�󯖯��)�;�M�_�
�*z�oomr�ZOOMIN�q��ؿ� ��� �ÿD�V�h�z� ��/ϰ���������Z*maxres��?MAXRES��	� ��p߂ߔߦ߸�[��� �� ��$���H�Z�l� ~��;ߡ����3��� � �2�D�V���z��� ������e�����
 .��;Q_���� ����*< N`����� w��/o8/J/\/ n/�/#/�/�/�/�/�/ �/?"?4?F?X?/i? w?�?�/�?�?�?�?O O�?BOTOfOxO�O-O �O�O�O�O�O�?__ '_�Ob_t_�_�_�_M_ �_�_�_oo(o�_Lo ^opo�o�o7a