��   v��A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����UI_CON�FIG_T  �x L$NUM�_MENUS � 9* NECT�CRECOVER�>CCOLOR_�CRR:EXTS�TAT��$TO�P>_IDXCMEM_LIMIR�$DBGLVL��POPUP_M�ASK�zA � $DUMMY�73�ODE�
4�CFOCA �5VCPS)C��g �HAN� � T�IMEOU�PI�PESIZE ޡ MWIN�PA�NEMAP�  �� � FAVB ?�� 
$HL�_�DIQ?� qEgLEMZ�UR� �l� Ss�$H�MI�RO+\~W ADONLY� }�TOUCH��PROOMMO�#?$�ALAR�< �FILVEW�	ENB=%%�fC 1"USER�:)FCTN:)WI��� I* _ED��l"V!_TITL�� 1"COOR{DF<#LOCK6%��$F%�!b"EBF�OR�? �"e&
�"�%�!BA�!j �Ơ!BG�#�!hIN=SR$IO}7�PM�X_PKT�?$IHELP�� ME�#BLNK�C=ENAB�!? SIPMANUA�pL4"="�BEEY�?$�=&q!EDy#�M0IP0q!�JWD8�D7�DSB�� �GTB9I�:J�<S�TYf2$Iv!_8Gv!k FKE�F�HTML�_N;AM�#DIMC4:1>]ABRIGH83s oDJ7CH92%!FEL0T_DEVICg1�&USTO_@ � t @A�R$@PIDD�BC��D*PAG� ?xhA�B�ISCREu�EF���GN�@�$FLAG�@ � &�1  h �	$PWD_ACGCES� MA�8��hS:1�%)$L�ABE� $T�z jHP�3�R�	� &USRVI| 1  < `��R*�R��QPRIƍm� t1�PTR�IP�"m�$$C�LASP ��)�a��R��R `\ �SI�	g�  �aIR�Ts1	o`'2 L1���L1���R	 �,��?����a1`�b�d~a�����y`� y�o��
 ��a��o�o1CU  �oz�����c �
��.�@�R��v� ��������Џ�q�� �*�<�N�`���� ����̟ޟm���&� 8�J�\�n��������� ȯگ�{��"�4�F� X�j���������Ŀֿ����`TPTX�����/�`� sȄ�$/�softpart�/genlink�?help=/m�d/tpmenu.dg���ϨϺ��� ������&�8�J��� n߀ߒߤ߶���W��� ���"�4�F�X���|��������������a�f�b�b�� ($p�-����T�?�x���a�a��c���c����l���c�R�ah�ah�h��2�h�	f���������`���`�  ���f ep���h#h�F�d��g�Xc�B 1~)hR \ �_� REG VED]����wholemo�d.htm�	si�ngl	dou�b trip�8brows Q�����u� ��//@/����dev.slh�/3� 1�,	t�/ _�/;/i/??/?�/�S?e?w?�?�?�?� H`�?�? OO$O6O HOZOlO~O�F2P�?�O �O�O�O�O_�E�	�? �?;_M___q_�_�_�_ �_�_�_�_oo%o7o Io[omooM'�o�o�o �o�o�o+=O as������ ���?>�P�b�t��� ������Ώ���O�� ���L�^�_'_��� ����ş�����6� 1�C�U�~�y�����Ư ��ӯ�o���-�?� Q�c�u���������Ͽ ����)�;�M�_� -��ϬϾ�������� �*�<�7�`�r�A�S� �ߺ�q���i����� !�J�E�W�i���� ����������"��/� ��O�I�w��������� ������+=O as������� ,>Pbt� ��߼���// �����^/Y/k/}/�/ �/�/�/�/�/�/?6? 1?C?U?~?y?�?Y��? �?�?�?�?	OO-O?O QOcOuO�O�O�O�O�O �O�O__�R_d_v_ �_�_�_�_�_�_�_��o*o�_o`oro�j��$UI_TOPMENU 1K`��aR 
�d�a*Q)*d?efault5_]�*level�0 * [	 ��o�0�o'rtpio[23]�8tpst[1[x�)w9�o	�=h�58E01_l.�png��6me�nu5�y�p�13�z��z	�4���q��]���������̏ ޏ)Rr���+�=�O��a���prim=��page,1422,1h�����ş ן����1�C�U��g���|�class,5p�����ɯۯ4�����13��*��<�N�`�r���|�53������ҿ�����|�8��1�C�U�g� y����ϯ���������"Y�`�a�o/��m!�`�q�Y��avtyl}<Tfqmf[0nl�}	��c[164[w��59[x�qG�y��tC8�|�29��o� %�1���{��m��!� ����0�B���f�x����������o���80 ��'9K~���2P�����\ ��'9K�� ����������1��/$/6/H/Z/U��|�ainedi�'ߑ/�/�/�/�/P��config=s�ingle&|�wintp���/$?6? H?Z?!Z�a�h?�?�e �?���?�?�?OO +O=OOO�?[O�O�O�O �O�O�O�O_a�%_L_ ^_p_�_�_�_U��_�_ �_ oo$o�_HoZolo ~o�o�o1o�o�o�o�o  2�oVhz� ��?���
�� .��@�d�v������� ��M�����*�<� ˏ`�r���������^��;�M�sc���;���s�� �}���e�au��X��@�F7L� ��`��t꒯4�j�X�6e�u7�����ｿ�Ͽ������27 ��G�Y�k�}Ϗ��0Ās���������!�1�M�_�q߃ߕ� T������������ 7�I�[�m����� ���������!�����6(�]�o��������$��746������)t<ϯ\�5	TP?TX[209©|Dw24§J��
�w18��� ���
�02��A#��[	�tv`�RxL.�u10�1����5S:�$treev�iew3��3��&�dual=o'8?1,26,4�O/ a/s/2�/�/�/�/�/ �/�/?'?9?K?]?o?��;/&�3$/6$�� �?�?�?
?#O5OGOYO kO}O�?�? "2�?8"�2K��O�O_�O��1��?�E��g_y_�_�6<_��edit��>_ P_�_�_o��/���_ �Cooo�o�oB�o�o ��oA�o�+ =Oas��o�� �����(�9��� Q�x���������ҏO ����,�>�P�ߏt� ��������Ο]���� �(�:�L�^�ퟂ��� ����ʯܯk� ��$� 6�H�Z��l������� ƿؿ�y�� �2�D� V�h����Ϟϰ����� �ϕo�o��o@ߧE� c�u߇ߙ߽߬����� O����)�<�M�_�q� ���W��������� &�8���\�n������� ��E�������"4 ��Xj|���� S��0B� fx����O� �//,/>/P/�t/ �/�/�/�/�/]/�/? ?(?:?L?��߂?1� �?���?�?�?�?O $O5OGO�?SO}O�O�O �O�O�O�O�O��2_D_ V_h_z_�_�_�/�_�_ �_�_
oo�_@oRodo vo�o�o)o�o�o�o�o *�oN`r� ��7����� &��J�\�n������� ��E�ڏ����"�4� ÏX�j�|�������a? s?蟗?�sO_/�A� S�e�w���������� �����,�=�O�a� #_������ο��=� �(�:�L�^�pς�� �ϸ������� ߏ�$� 6�H�Z�l�~�ߐߴ� ����������2�D� V�h�z�������� ����
����@�R�d� v�����)����������ƚԔ*de�fault%��*level8��ٯw���? tpst[1]�	��y�tpioG[23���u����J\men�u7_l.png�_|13��5Ж{�y4�u6 ���//'/9/K/]/ ���/�/�/�/�/�/j/ �/?#?5?G?Y?k?�"�prim=|p�age,74,1�p?�?�?�?�?�?�"��6class,13�?*O<ONO`OrOOB5xO�O�O�O�O�O�#L�O0_B_T_f_x_{?�218�?�_�_ �_�_�__B6o9o�Ko]ooo�o`�$U�I_USERVI�EW 1֑֑�R 
����o��o�o[m �o'9K] � ����l��� #�5��oB�T�f���� ��ŏ׏鏌���1� C�U�g�
��������� ӟ~�����v�?�Q� c�u���*�����ϯ� 󯖯�)�;�M�_�
��*zoomr�?ZOOMIN�q� �ؿ���� �ÿD� V�h�zό�/ϰ����������Z*maxr�es��MAXRES��	ߧ�p߂ߔߦ� ��[����� ��$��� H�Z�l�~��;ߡ�� ��3���� �2�D�V� ��z���������e��� ��
.��;Q_ �������� *<N`�� ���w��/o 8/J/\/n/�/#/�/�/ �/�/�/�/?"?4?F? X?/i?w?�?�/�?�? �?�?OO�?BOTOfO xO�O-O�O�O�O�O�O �?__'_�Ob_t_�_ �_�_M_�_�_�_oo (o�_Lo^opo�o�o7a