��   ��A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ������DMR_S�HFERR_T �  $O�FFSET  � 	  /GR�P:� $�MA��R_DON�E  $OT�_MINUSJ � 	sPLzdC�OUNJ$REF,j�PO{���I$BCKLSH�_SIG�EA�CHMSTj�SsPC�
�MOVn �~ADAPT_I�NERJ FR�ICCOL_Pz,MGRAV��� HISID�SPk�HIFT�_7 O �N\m�MCH� S��ARM_PARA�O dcANG�o y2�CLD�E7�CALIB�Dn$GEA�R�2� RING,��<$]_d��REL3� 1� N �CLo:o � �AX{ � $PS_�T�I���TIME� �J� _CMYD��"FB�VA >�&CL_OV�� oFRMZ�$DE�DX�$NA� =%�CURL�qW���TCK�%��FMSV>�M_LIF	���'83:c$�-9_09:_��=�%3d6W�� �"�PCCOM,��FB� M�0�oMAL_�ECI��P:!o"DTY�kR_|"�5:#�1E�ND�4��o1� l5M�P P�L� W � � $STA:#TRQ#_M��� KNiF�S� uHYsJ� hGIʀJI�JI�E#3ApZCaB�A� �$��ASS> �����A�����@VE�RSI� �G�  �QIRTUAL�OQS� 1X +���N ��x_ c_�_�_�_�_�_�_�_ ofP��6me Q^o�Lm���=�����a�� �?_&���#Ko�o Goql�o�o�o$�kW]rF������d�������=L���8�?�9���@�Y�~����� ��Ə؏���� �2�D�� 1Uo�}�g����D  2�Ο�� ���(�:�L�^�p���<��������Я� ����*�<�N�`���2P��(�������� ܿǿ ����6�!�ZπE�~�iϢύϲ�����$4 1N\����H��}Id��J$�F�5�WSPN�K"[�!��IC߳H���FGʛ2P�(�>x:C���A��]߶τ� �߁ߺ�U�gߡ��߀��1��U�@�y����V�aV�q"t���� ��� p���l����1�C����%��345678901c�k���� ������������`� "4��
��d��� v����J� *N<r��� ��\�//8/ ��q/���/"/�/ �/�/�/T/%?7?�/�/ j?X?�?|?�?�??�? >?P?�?�?OTOBOxO �?�?�OOO�ObO_ �O_>_�Oe_w_�O,_ �_�_�_�_�_oZ_+o ~_�_
o�_^o�o�o�o o o�oDoVo$�oH 6X~�o��
l ����2�D��k� ��J����ԏ�� N�`�1�����d�⏈� v���������J��� *��N�<�r���ڟ�� �����\�ޯ��8� ����q�į֯��"�ȿ ��ؿ��T�%�7ϊ�� j�Xώ�|ϲ������ >�P��Ϝ��T�B�x���ۙ��ϱ��,���8����U��$PL�CL_GRP 1�o�� {p(�?�  "� 4�,�W�(�{�f��� �����������A� (�2�t�