��   g�A��*SYST�EM*��V9.1�0214 8/�21/2020 A   ����BIN_CF�G_TX 	$�ENTRIES � $Q0FP�?NG1F1O2�F2OPz ?CN�ETG  �DHCP_CTRL. � 0 7 A�BLE? $IP�US�RETRA�T�$SETH�OST��NSS�* 8�D�FACE_NUM? �$DBG_LE�VEL�OM_N�AM� !� FTޒ @� LOsG_8	,CMO>�$DNLD_F�ILTER�SUBDIRCAPC�  D��8 .� 4� H{AD_DRTYP�H �NGTH����z +LSq D� $ROBOTyIG �PEER�ބ MASK�MR�U~OMGDEV������PIN�FO�  =$$$TI� ��RCM+�T A$( /�Q�SIZ�!S� T�ATUS_%$MAILSERV� $PLAN� �<$LIN<$�CLU��<$T�O�P$CC�&F�R�&YJEC|!�Z%ENB � A�LAR:!B�TP�,�#,V8 S���$VAR�)M�O�N�&���&APPL��&PA� �%��'P�OR�Y#_�!�"A�LERT�&i2UR�L }Z3AT�TAC��0ERR�_THROU3US0�9H!�8� CH- c%�4MAX?WS_�|1��1MOD��1I�  �1o }(�1PWD  � cLA��0�ND�1�TRYFDELA�-C�0G'AERSI���1Q'ROBICL�K_HM 0Q'� XM�L+ 3SGFRM2U3T� !OUU3 3G_�-COP1�F�33�AQ'C[2�%�B_AU�� 9 R�!�UPDb&PCOU�{!�CFO 2 
$V*W�@c%�ACC_HYQSNA��UMMY1oW2�"$DM*� $�DIS�� SM	 l5�o!B�"%Q7�IZP�%� ��VR�0�UP� _wDLVSPAR!#R�PN,#
3 �_��R!_WI�CTZ�_INDE�3^`O�FF� ~URmiD��)c�   �t Z!`MON��cD��bHOUU#E%A�f�a�f�a�f�LOCA� #$�NS0H_HE����@I�/  d�8`ARPH&�_IPF�W_* O�F``QFAsD90��VHO_� 5R42PySWq?�TEL�G P����90WORAXQEF� LV�[R2��ICE��p� �$cs   �q��%
��
�p�PS�A�w�  �5�	�Iz0AL��X' �
���F���P��!�p�i��$.� 2Q������������ Q���!��q����$� _F�LTR  �\�� �����������$Q�2��7rS�H`D 1Q�" P㏙�f���ş ��韬��П1���=� �f���N���r�ӯ�� �����ޯ�Q��u� 8���\�������󿶿 �ڿ;���_�"�Xϕ� �Ϲ�|��Ϡ����� ��6�[���Bߣ�f� �ߊ��߮���!���E� �i�,��P�b���� ������/���(�e��T���L�����z _L�UA1�x!1E.��0��p���1��>p�255.0��&r��n���2����@d %7I[3e���� ����[4 ���T'9[5U���{���[6���D �//�)/s��QȁM�A¸MA�H������ 'Q� ��u.<�/? &?�/J?\?n?A?�?�?m�P�?�?�?�?�?O .O@OROOvO�O�Ou.�kOl�q��O�L
�ZDT StatusZO�O5_G_Y_n��}iRConn�ect: irc�{T//alert ^�_�_�_�_mW#_o@o,o>oPobot�^�d~2g���go�o�o �o�o�o�o	-?�Qcul�$$c9�62b37a-1�ac0-eb2a�-f1c7-8c�6eb57836fe  (�_�_ ���"�p�1!W��(��"S��JE�� 0X��C� ��,$��� W���ˏ���֏�� %��I�0�m��f��� ��ǟ�������!���u�R����� D�M_�!����S�MTP_CTRLg 	����%� ���DF���ۯt�ʯ���'��Lz�N��!
�j��y�q�u�����Ԙ��#L�US?TOM j�������  ���$T�CPIPd�j���H�%�"�EL������!���H!T�P��j�rj3�_tp�b;���i�!KCLG�L�i�|��5�!CRT�������"u�!C�ONS��M�[�i?b_smon����