��  	c4�A��*SYST�EM*��V9.1�0214 8/�21/2020 A  �����AAVM_W�RK_T  �� $EXPO�SURE  �$CAMCLBD�AT@ $PS�_TRGVT���$X aHZ�gDISfWgP�gRgLENS_�CENT_X�Y�gyORf   �$CMP_GC}_�UTNUMA�PRE_MAST�_C� 	�G�RV_M{$N�EW��	STA�T_RUNARE�S_ER�VTC)P6� aTC312:dXSM�&�&�#END!OoRGBK!SM���3!UPD���ABS; � P/ �  $PA{RA�  ����AIO_CNV�� l� RAC��LO�MOD_wTYP@FIR��HAL�>#IN_;OU�FAC� g�INTERCEP6fBI�IZ@!�LRM_RECO�"  � ALM��"ENB���&O�N�!� MDG/� 0 $DEB�UG1A�"d�$3�AO� ."��!_I�F� � 
$_ENABL@C#T� P dC#U5K�!CMA�B �"�
� �OG�f 0CUR�R_D1P $Q3LI�N@S1I4$C$AU�SOd�APPI�NFOEQ/ 9�L A ?1�5�/ H �7�9EQUIP �2�0NAM� ���2_OVR�?$VERSI� �� PCOUPLE�,   $�!PPV1CES C G�1�!�PR0�2	� � $SOF�T�T_IDBTOTAL_EQ� �Q1]@NO`BU SPI_INDE]�uEXBSCREE�N_�4BSIG��0O%KW@PK�_FI0	$�THKY�GPAN�EhD � DUMMY1d�D�!U}4 Q �ARG1�R�
 � $TIT1d ��� �7Td7T� 7TP7T5�5V65V75V85V95W05W>W�A7URWQT7UfW1pW1zW1�W�1�W 6P!SBN�_CF�!�0�$!J� ; 
2�1_�CMNT�$F�LAGS]�CH�E"$Nb_OP�T�3�(CELL�SETUP � `�0HO�0 P�RZ1%{cMACR=O�bREPR�hD0�D+t@��b{�eH-M MN�B
1��UTOB U��0 9DE7VIC4STI�0�A� P@13��`BQd�f"VAL�#ISP�_UNI�#p_D�Ov7IyFR_F �@K%D13�;A�c��C_WA?t�a�zO�FF_@N�DEL�xLF0q�A�qr�?q�p�C?��`�A�E�C#�s�ATyB�t�d�MO� ��sE � [Mp�s��2�REV�gBILF��1XI� ~%�R  � �OD}`j�$NO`M�+��b�x�/�"u�� ��Ԯ�QX�@Dd �p E RD_E�b��$FSSB��&W`KBD_SEV2uAG� G�2 "!_��B�� V�t:5�`ׁQC �a_ED|u � � C2���`S�p�4%$<l �t$OP�@QB9�qy�_OK���0, P_C� y��dh��U �`LACI�!��a���� FqCOM9M� �0$D��ϑ��@�pX��ORB�IG�ALLOW� �(KD2�2�@VA�R5�d!�AB e`BL8[@S � ,KJq�M�H`S�pZ@M_Ox]z���CFd7 X�0GR@�z�M�NFLI�<��;@UIRE�84<�"� SWIT=$/0k_No`S�"CFd0�M� �#PEED��!�%`����p3`J3tV�&$E��..p`L��ELBOF� �m��m��p/0��CP�� F��B����1��r@1J�1E_y_T>!@Բ�`��g���G�� �0WARN�Mxp�d�%`�V`N�ST� COR-�rFLTR�TR�AT T�`� $ACCqM�� R�r$ORI�.&ӧ�RT�SFg C�HGV0I�p�T���PA�I{�T��P��� � ��#@a���HDR�B��2�BJ; �CѪ�3�4�5�6*�7�8�9�4���x@�2 @� TRQ��$%f��ր�׍��_U���ѡ�Oc <� �����Ȩ3�2��LLEC�M�-�MULTI�V4�"$��A
2q�CH�ILD>�
1��z@T}_1b  4� STY2�b4�=@�1)24����=�� |9$��T�A�aI`�E��eTO��:�E��EXT����p���B��22�0>��@��1b.'���}!�A�K�   �"K�/%�a��R���?s!>�O�!M��;A��◒M�� 	�  8=�I�" L�0[��� R�pA��$J�OBB������TR;IGI�# dӀ�� ��R�-'r��A�ҧ��_M��b$ tfӀFL6�BNG�A��TBA� ϑ�!� �
/1�À�0���R0��P/p ����%�|��Bq@W�
2MJW�_RH�CZQJZ�_zJ?�D/5C�	�ӧ��@����}Rd&� �����ǯ�rGӨg@NHwANC��$LG/���a2qӐ� ـ@��A�p� ���aR��>$�x��?#DB�?#RA�c?#AZt@�(.�8����`FCT����c_F࠳`�SM��!I�+lA�%` �`  ���$/�/����[�a��M�0\��`��6أHK��AEs@͐T�!�"W��N� S'��I��'  �. II��2�(p�STD_C�t�1Q��WUSTڒU�)#�j0U[�%?IO1���� _Up�q�*c \��=�AORzs Bp;�]��`O6  RSY�G�0�q>EUp���H`G�� {@]�DB�PXWORK�+~* $SKP_�p���DB�TR�p , �=�`����Z m�OD3��a _�C"�;b�C� �GPL :c�a�tőS�D��G�Bb����P�6.� )DB�!��-|B APR��
���DJa3��. p/�u����� �LUYI/b_����0�_^���PC�1�_�tS~�EG�]� 2��_�S6PRE.��R3�H $C��7.$Lc/$USނ�z )kINE�7A_D1%�ROyp��ŀ����qbc7 T@zfP�A���RETUR�Nxb�MMR"U���I�CRG`EWM��0�SIGNZ�A� ���e� 0{$P'�1$P� &m�2�`��`tm�pDIp �'�Bd.a|	r�GO_AW ����0ؑB1I�CYSd�(�CYI�4��B�`1wsqu�|t2vz2�vN�}��E]s�DEVIS` 5� P $��RB���I�wPk��vIG_BY���p�TQ޻tHNDG�Q6� H4��1�w��$DSBLC��O��v�G@��SP_qL��70/�F@]�d�FB���FERa8����t]s��
�8> i�T1?���MCS솀�FD ���
[2H� W��EE���p%F��ŻtSLAd��09  ��INP�^��]�`�]q��:P +8�S��0x�`^���^���FI�2�������A	A9Wl���NTV�㜒�V~���SKI�#T�E����a���T1J�_�#;2_�PD�SA�F�T�_SV�EOXCLU�῰�%D6@Ll �Yք��3�HI_V
0\2PPLY�@0«�G������_ML%��pVORFY_�C��M��gIOC�UC_� ����O�p��LS(�`M2&T4�A1��s	���@PdE&�gp�AU��NFK6u��upZ��pm�ACHD��O���^���AFC C	Pl��TD�4P~�� N�� ;�P@T�ќ�0,@ �B��N���=� <Y���TĲ�?� ���{�SG5N��=;
$�` �a>aR0I�3�g@ _B�M�_B]�ANNUN��P~��ÅuC.@ �`/�ɢ�� �����2�EFC@I�R>p�c$F���4OT�` {�&TD�(RQ<�#QI�-Mb�NI�R?��4��6�A��R�DAYCLOADz�T-��'S5#Q�EFF�_AXI��@�P�QO3O�йS�@_RwTRQ��A D1�t	`��Q,@ ��!EVp�Ӓ���@�0}��0��{��MP�E{� BV������$s��DU�`���.�BCAB��C���P�NS"�+0ID�W�R���V!� V�wVq_���V �DI� ��4D� 1$V�`SEm�TQj�}�'���D�^E_ln�$�VE� � SW���[a���2��A��OH��)�3PP��%�IR�1Bu@p�&���b���� ]�w3W�O � W��vM����C�0��cp��RQ�DWF�MSw0��A�X,���$�LIFE �@����-Q��N�������Co���CB0LqN]a�f��OV0HEQ�NSUP�K2��"�@_oS�1_��Gq�Z�
W�
B1�0�#��@�k2XZ_ LQVY2�C9`T_@D``��N�����J�! >�_� ��F� �4�E `�pCACqH,�\�]SIZ(�T ���bN�UFFI� ���@(T$��'S6.ҍAMp0��F 8��KEYI7MAG�cTM,aV#���a�^�hB1�OC'VIE�aG�2� �L��H���?� 	R��D� PH���ST'�!C"D�K$�PK$��K$��K EMAILK�u`[��0��/FAUL�RI�2sc�C� COU�0iA�0�T`�1J< �$�#�S�m�ITW�BUFp��p�t��0�0n B�$�tCු���"�3� SAV -5�"����H7@@���P44�
`�N�_0� 5LЉ9OTgb+����P�P�:���7AXC����X� T�a3�_G��
��YN_\N� K <\�D�uTPb�M�M8�H 5TL�F~`$�`��DIزE�@`�aILY���G1��&G��Da:AF����baMa�`A�#�3C_^`��`Knd�@^DQ�Rp��E�(ADSP�6BPC�KIM:3�C�A��A��U�Gd meڠ� IP��C7�3��DTH���B��T�aa�CHSEC�CBSC	�"�PV���Z�P��3�Tp��NVk�G �S�T�F� F���0ad�C5@�1aSC���u�CMER��QF�BCMP��~@ETn;� N�FU� �DU� ́�`���CaD�IYP�0�# ��`SNOu�=�O���p�zbL�xds�P�zbC""��e
��2�!uc|�0� PH *�aL��_c�q�1f��,� '��dD��f"��f���fP���f��f7�i8�i�9�j���hz1z1�z1(z15z1Bz1�Oz1\z1iz2wz2T{z2z2(z25zU2Bz2Oz2\z2iz�3wz3z3{z3�(z35z3Bz3Oz3�\z3iz4wr �EX	T��=�QB\h@%�@�e@C��e�0F{DR��RT� �VW��2�򁑇R��R�EM��Fq��OV�M�C��A��TRO�V��DT80КMX�ߜIN��: Ϛ��IND���
�F@�0@G�1d�ِ9 ��9D��ِRIV԰&���GEAR�AIO��K��$�N5@���������� %�Z_MsCM� ���Fe ;UR3bS ,�a1�? 9 P?\���?�E,� �� �1`v�T0Ч�5P�1��RI^eJ���#ETUP2_ gU ���#TDGP0��$Ti��Z�T�qa��"BACBV T(D��"eD)_J%�ýc0@ѰIFI:�0@`��`�Ь�PT�����FLUI6$�W �� (� UR t�1@�2MA�P� ����I��$(�Sܰk?x4�Jb@CO|0Ο3VRT$���x$�SHO�ѱ��#AS�SjP�1(IPQ�BG_����s��s��(s<��5sFORC�"7�^�DATA��X�"KFUס1:B��2:A�LOG���Y �|*�NAV�0)�(�X����S�"&?$VISI[��SC�4SE�t�7�UVB�Or���Bòx�A�Z�$PO,��IE��FMR}2s�Z �� i`f⁑s@�օ��������ǖ� �堒_wqX���IT_ֱSd���ME�j�|�DGCL�F;�DGDYd�L	D�H�5
?�ѡ�Mcp8#[���� T�FS�07$\� P2���sC�0$GEX_������1�0��PE��3�5��9G�Q��] ��0b�SW5O��DEBcUG��]�GRc���U�SBKU`O�1�p  PO@�Ј�t�"`G�t�Ms�gLOO�3��SM��E<2qa�& _E �^ �j��T�ERM��_���!O�RISA��`��cp�GSM_`@]���a������� b��~�UP>"c� -�D�^(���f _>�G�k
}�ELTO�!>B�PFIGf?Aנ�S�`b`$UFRfB${`�� �Ne�OT��PTA�iP���NSTT@P�AT^Qi�PTH	J&aL`E9 d2U`�ARTU0�� U1�"�>ARELAc1SHCFTPR?A3__�QR/`Ic ) $8��b.႐S�S�2SSHId+�U�b O1AYLO.P�1 A���j����e[PERV p�$��T@�A��Ȱ+%��ȰRC<��eASYM3A�eF?AWJ�$� �E$�/[)�OaU$T@ A3��&IPS��Q֯ORT@M��/����d��t���� �1)`HOs���e� �˶s�i`OC���$OaP^��A�cv���$a�i@��R0R�S"�OU�Se�R��5m8K��e$P�WR]�IM�5"R�_H3(*� ?AUD$�kSVoc1SD]fH�$HdE!@�ADDRC�H��GP7A,A%A�t`RE�.�ag H2�S�PFр��dE��dEsdE(sS�E��H��`HSY`MN�hW�@0��"QebaOL/SW�{0xR�\f��ACRO��<��ND_C/Szbx��4�QROUP�SB2_��
Ғ�11�q ��:S�DY3 DY��EX@pDY(pDY����AC�<��SAVED?W�S�OUG�C��i $��@0_D)���j«B�PRM_
�~�H�TTP_z`H�aj; (;`OBJB�%B6��$C�LE�0|a�`k � 4���6�_�T��XbS�0�3��KRL�9HITCOU����G�LS�j0Xbb�$�f�j0�ʷk0SS���dJQ�UERY_FLA��C_ _WEBSOCI��HWcq�+��l_@� INCP	U�R*�Ovma��K��0pzD/q�D/qǂ��IOLN��m 8�2�R��i�$SL���$INPUTM_��$�0~xPy�7  ZpSL�P+�nep{�u�tB#�u�B"NAIO�PF_A5S��o��$��B�
�qN�Y��2��0ksM�ts�HYB�5����A�pUOP��p `�pS�C���%���,�}��0P�3�0s����,������IP_M�E\��q X�pI1P,@�Rւ_NP��`*�G2B��O��B�SP���P���BGȬQ�-�M<!�r �l �TA�3`As�TI���%� ��_��OPS^�BU��I�D�Ўbs���x0�� c�
,���� s�r"?�r�S��pNҘ���ӕ�IRCA_C}N� t �Jim�pCY�@EA� �C��q��31�#��@xz"���!DAY_����NTVA����u�p�r#��u�SCA�Fu�CLO᎑j����@��u��ڔ$��N_R0Cβ򐎒c�6�v�r��^3%���'b������Pi��� 2�u �p.����wp��\�'b\�LAB��z��Ѐ�UNIбn�	 ITYl�.�0E"L�R; G���x�r��R_URLЀ$A�AEN|�k�*��0��CT�AT_U#� ��Jp��yр$�_%E�pRk�.���AS��q8�J�aC�F�L��K��P
W�r�
��UJR�%z ��J`F��(����D�£$J7S%�J�8��7&�h�����7����8�ɭ�APHMI�Q����D���J7J8"�L_�KE��  ��KQpLMܑ { <٠XR�p$p��WATCH_VA��A�ű#fFIEL��"Cy�2Ҳ�| �
��V�G-1��CTpܰ��� �LGɳ�}� !�LG_SIZRdv��հ�����p��FD��I ���ة����������� d3��V��V��pV��@V���V�K!G�� _� _CM�������AF�!�����А4(������������p��� �I��
���0��������RSU�o  (��LN��j�"~_��`DE��E�r!�s���S��0�L���DAU��E�A�PQp44���GH�52X��pBOOYA�� C�ʀIaT�c��� �RE4��SCR��|c�D��PKr,QMARGI �q�;�v�S4e�d�qS8c�rWC�q����JGM�MNC�H���qFN(ҞK����	UF����FWD�HLSTP�
V�������RS?H� ��C�~"�� w�U�Q�v����2�G�	PPO�"�2�� ��	EX.�TUI�I;�� �;�8bZ#�Z#� ����R��P# #N�A�3ANA�rA1���AI���D�� �DCASf�lC�#zC�"O�(EO�'SK�2�(S�(ZIGN�Ў������4��$DEA|LAL"�Xp�q���Ѐ����T��$�׳�rh
���AA��С۠lp*s�A��S1�52�53�1��"� �Ђ �Jk�0�$�u�t���Q�e�X��:FSTe�R���Y�B\A �$EkFCkK���PzF�F8{�$�у Lp#� n�8����Co`��d�P��D�5#_ � ��Pt��P��$ Sm��MCt�� ��J`CLDPe� �TRQLI��"�PY>T�FL%�iR�QrS��D��rWpLDrU\TrU�ORG(�v�R��RESERV2t�T>s��TIr�/Sv�� �� 	[UvMTrUS�Vd�PP^�	�Q+d>3fRCLMCAd�_��_SiTp3al0MDB�G�qͰ�?�$DEBUGMAS&�(_�P���UuT� |��E�����MF�RQV�� � ���HRS_RU��q�A'�A5��FgREQ����$� ��OVERt���tF��P�EFI��%�A(��a��b�Tǉ \�q��$9U@%�?`��SPS�0C�	sC��BcN��sScUݐ�a�?( 	��MIS�CuŊ d}�AR5QA�	�TBN ��c �m!�AX ��-��.�EXCESH�{��rM��̱���a�r Ŀ��rSC@� � H"�	�_�S��8���,�>�.PK�ɴ��r��N �eB_^��FLIC�DB �QUIRE�MO���O�pv�QL�@Mȵ� P��E���4�Ab�aND��q�Bހ�{�r��؄�D��>��INAUT4��GRSM����+0NfB�n�j�|�r�PST�Ḻ� 4٠LO�CFRI��EEX��ANG�"�q�aO[DA�e��p|����MF���Cv7I��BA �Eq�o�fSU�P�FxpFX;�IG}G � �` �Cn�(�C��Da�br \B��^@ɨ^@ئ���P��7�qTIvл�ypro�M+��b� t9�MD6���)D�� O��XaL�H���O�DIA��P�>�WiO��1�O�D��)/�t�)`nހ� m�CU�СV��#`�qՁO\_�`y�� ���CC�L�`rr�� �P �hJ���P��KE�^���-$B+p��@�ND2ZbZ�P�2_{TX�DXTRA�#4|�lb�E�LO��ހ1�k���� ��u��ǲ�ƪ�%�RR2>�u�� .�����A0a d$CA�LI�o�G�!��2��0RIN����<$R��SW0_d,�lcwABCJ�D_Jb�����pC�_J3W�
�Q�1SP�Т��pP�Q�x�3w�̱�@�pB��Jlc���R(aOu1�IMl`�rCSKP _Z�Ի��#��J���r�Q��������_cAZ/b��I�ELZ1<��ZaOCMP��q��q��RT�at��11��В��1���{ :��Z��SMGY'�vzdJGPSCLN�
�SPH_0�p7���㓰�p��RTEIR+���� ��_� 
)Q6@A\ SC�r'�sDI_���23U��kDF�0H�LWN�7VELPQIN�Bf q�_BL� �ry���³qJi�~�����MEcCH�2lbwqIN
�q���ǲ��]�q��:�@_�p �����/��0�􆂛��?�Հ�DHN�~�����0�$V������{!$���'q
�A�$O1�`R�����H �$BELZ��g��_ACCE� x�la� IRC_(��a�PNT�q;C�$PSN�CRL�0 ��XS���?�� � G��	�3�ؠQ�_�1lIO"u�pn�_MGsDDl(�
�FW3P(���ظ�}DE�PP�ABN�RO��EE_�1�PP��1�a�����0$USE�_���#P+pCTR��$Y�~ .a �AYN�pAm 6&��f�6!!M�aұ�"fOk�
c$INC�����p��'���ENC��L��r���� I�NCBI��%)���N�Ti��NT23_L�
��#LO]�
�09pI\��6R���p����0����C���&MOSIq��߰O!s��rPERCH  ��7q� y7��3� 2zd�o�g� %&N��AC�5L$�ӻ�����%��:F36TRK��AAY���3�� HACWELC�z暁�"�`MOM}"����P̰����cC����DU��DS_BCKLSH_CC �E�`X68p>#�s�C�"�ZM!�CLALM��$�a�@ 5UCHK����Z�GLRTY@��A��$��Q'�_f�NM4_UM�c�VC�cpz��SpLMTtЃ_Lj b�Tv��WE �]�P�[�P��U���0�c�2 d�8PC�1�8�H��&�p�UCMC���z~CN_	�N���f��SF��9V  "��'�TaC�eXh7CAT�^SHf�	� ~�&yQ�A�&�����̗�mPA�T�"_P�UrC_����OFm0��_CqtbUJGJ�d�es�W�OGrg�TORQU ��K3hI��0c2��r_W�EHD���m�t^�ud�uI*�{I
�IdF0��q���I���vVC� 0����j�1p�n��0�v�JRKp�������KDB��M����M���_DL^�2GRV��t�^�dՁH_p��Ӄ"�COS/�|�/�LN��R�s�Y� ^ T���T�&���~�D�bЅZM�c6ՁMY[��Θ;�I�C��THE{T0#5NK23d��X\�CB�CBXC��AS�C�&�0Q�^Q��SB^o�N)�GTS���C{��Kq��:s�祪��$DU_P�7ʢ��٧ʏ�Q�1_4cqNE
��KoT��-�< �A�:�C�!�,�,��LPH/���%�S s���~����������(����:�V\�VQ�N �t�V��V��V��V���V��VȻVֹH�\�u�{�s��a�Ȑ�H���H��H��HȻH*ֹOM�O\�O�r�UO��O��O��O��UO��OȻO��F��>���~���O�SPBALANCE_ޑ���LE��H_�S�P��o���~��ҍ�PFULC�����썕��1���UTOy_ZPbUT1T2^��2NAQ�� ~���@�A������AT	@�OA��pINSE9G�<1REV��<0��!DIF2E	1�l��?�1�%@OB��%Q���G2�p� LQ݄?LCHWAR�SABAq�E��<0ސ(U!���SXUAPdt�83�?S�� 
u��qܗ�%ROBm0CR�C��ib  �C��_]rT � �x $WEIGHR p$M���tp�IR!0IF
!�LAGC""bSC"��C"7BIL)OD�@?0&ST� P��%PB  | �`�������
� �D!]q  2y�J4DEBU�LXɠMMY�9���N+s�p3$D�1$� op� �   �D�O_� A�� <@��rh��D!0�BB�: N�#_!0D �_O2P ��� %�PT� �!�QTx��� TICK-�T1� %j�@s!Nm0M�	m0R�@D!�=�=�� PRO�MPR#E/� $IR�pB!hP��0"MAIڀ}!T"�_# ���^AV �R�CODwFUJ ID_�0'%������G_SUFF�&� 9!��DO����< �GR#=�e$�q$=�|%=�%�qe$�� ����H�_FIv�9�#ORDB ��36b�"B!� �$ZDT.%���_��4 *��L_NAs52>�DEF_IE852 �Q4�I�S�}3��5�IS��`���3�O4�a�4�abSDQ��B�4�wD�pO�� LOCKE+q_#����1e"_ UMd%52e$ }3e$�5e$�2q"gCp% `3q$�4q"Q�F�1|# H�^q|%52|%}3|#�GUa(8P�4H�1D�� WFHEU<Cxp��TE0Q��� LOMB_t_RzW0VIS=�WITYAoqOCA_FRIN�S�#SI�1�Q�Rp�W�{�W3�W�XW��[倩V��_i�!EAS�"�q�Tp@T��V4�Y5�Y6�ORMULA_I�+q�G%7� h� �7�COEFF_OW��dW���GqS �CaA���_GR�� � � $h<@��
XGTM/G�'t<E]DCA|ER���T%D$4� �  �G�LL�$@S/�_3SV�4�x$hV� q����d� � r�SETU�3MEA��D b� _�"��� � �p��  � �` �� �A�:2�sA0AD�b �Q�";��@�1@�G����RECt�!�2SK_���s� P��1_USERz��,�8����z�VEL>����,�����=�I0f���MT8CFG���O  u��Oc�NORE�� ���-��� 4 p�s^�d�XYZ�#�f������_ERR�� ��ep6 A�c\�}��Ҁ� BUFINDX1�t��PRt� H��CU\�d��1xӃ���!$������10�dQ���G�r� � $S�I�`�P �ᝀVOx
����OBJE��ADJU����AY9p���DJ�O�U� 5���C!�"=��T��y���x��DIR}��������⎴�DYNb�b��T�R�5�R�QHB 4���OPWOR� ��,� SYSB9U*�2�SOP��$�q�U���P<@߂4�PA���6�_�2�+OPz U4�(��xt�e�IMAGo�1��q�SIM���IN`\���RGO�VRD��%���g�P i��������@ C׵d��L:@BY��� �PMGC_E0��N*�M±�1�2��sSL���� ���OVSL��S:RD#EX�1�0K�2c���a_��cǬ ��cì  mÂ�}Ȫ��C��70����Ƿ�_ZER� �*��s��� @h"���~�O0RI���
��������T��'�L�����T`�W ATUS�p�C#_T����O�B+pYրB���3�.�0��� D�e�N�LҾ��`M��!��o��XES� ��һ҆��ò�����R�UP:��0�1PX��y�b��3ǂ���PG텳��$SUBA�~��AA��JMPWAIT��r�Y�LOW/�^�' CVF�vc�\�R���q�CC��R���i��IGNR_{PL�DBTBW P�1d�BW ����U*��IGL��I�c�TNLN����R�֡5B�PN�E�PE�ED��T�HADO!WW b���ES�M��b�+�P0SPD��� L��Ar�Q0m�/��{�UN �y���R�м�LY0��K��_PH_PK����?RETRIE��bi�'����FI�Ƕ �:����� �2���DBGLV~��LOGSIZ���1KTy�U�s2D�8� �_TX�EMB�`Cn�F�X ARR|.R+�CHECK��N1��P��p�c������LE�4pP�A#@T��C�O��P4��p�bAR%"���#�1'�O� 0��`ATT���x�%X 0��1��UX�����PL,  $���/QSWITCH�T��aW�AS����SLLBp��� $BAv�D
C2�BAM�������J5L����6�|_KNOWh����U=�AD���`x�D��)PAYGLOA��@%#_���.'�.'Z+#L�AA��q�0LCL_ʐ !�pg"�Ӂt$*˲�&F�)Cgpb*(�e$�`Ib(Ripb'${�~$B7`ʑJE��!�_Jl!��֑ANDz�U�
4l"�!(�"a�PL�AL_ ��`x�ѐ����PC�>�D*#E=��J3�036� T�`PDcCK�22�CO�p�_ALPHC3�3BaEБsaC?U< ��b|��� � �.�$/D_1+*2U$D�pAR��H�5FC^�TIA41I51I6>�MOM��=C]C�JC]CWC�Bp�AD�=C�FJC�FWCPUB�RbD�EJC�EWB'��@30ʑq�  �� MO"L� ��T���� e$PI����3��0'P&Y��J)&YI2[I@[INS�DS�V�V�ޠ2������1�HIGo1�q�j��Vj� q�����V�S�X���Y<��q�SAMP�Я��:d�W;cq�3 �piaʐS�Œxd� �fj��0�i@Œߠ䢐:@�e/0��H��cIN�l/0c�h�k�dq���jx�d{2{GAM�M�eSU�A�$G#ET�R��3�D�4҂;
$60IBR���]IL�$HI:�_��H��Œ�vEѐ�xA�~�p�vLW�}�v�|�y@��v�2�V�51C��GCHKİ��q�x>I_`�ޔ.2�8.1��e|�uCޔ�F{�33 ��$e8 1���I�RCH_5D����RNs�8���LE���R����8�Ѐ��MSWFLܡ��ASCR�100{�. xd39]��g�ʐ=@�iq�j���PI�3AVMETHO��æ��妒AX$���X4�p�ERI���:d3fsR�� 5	D�Q�0FWt;ac��c�(�L�;a=�OOPa֑S��a֑'APP��F� 0W�x�c��cRT��2�O0j�0�������DR 1�%��D��ѪNP�ѢRA� MG�vOSV	Q�P; �CURC��GRO<7���S_SA�ܴ,5���NO�0C���� �45��t�?6/H/TX�����zP��UϸCDOi�A�rdyes��e�X ��W��X3�/��k#����D�T� � ���YL$S�!�g���S�"6A9��K����!�����!_�C����M_Wd���C�����?�M���ˇ ��21~�L�T�K��r PM&�R� ��}�R��WE�S$��L3X!EШ4Cү4@CҶ4C�W4���pN�P�sf��/0X��O�3�.1Z�� P{�T� ���M��z�w����������4@������L:�1_Z� |v1�� 5�]I��JC��WC5�6J ���PJuuMs���ſ�Y s�P��PMON_QU?`� � 8� QCsOU��QTH_�sHO~�:�HYS3ES�:�UE%�+��� OX�  ��P�#ПuV�RUN_T�O���g�R
P� P! ��C�����INDE�ROG�RA��J��2C�N�E_NO���ITx�A��g�INFO��� b������u��I��� (SLEQ�V"�U" ̺�A�OSU���{ 4� ENABq�>��PTION
�ERVE�R~�Q��VGCF_� @b.�J �.1����p�R��m��@EwDIT��� �R�R��K�A�S�qE�psNUAUTQ�	COPY�A�P*�Q]�M�qN48M��PRUTR ;N� OUC�Q$G���?�RGADJn��� hv0X_��AI���п�пW��P����S��rN^0_CYCq��/RGNS[�s�=��LGOZ��PNYQ__FREQ�BW�`��VP!SIZn[�L�AœG!�XC�`�UCcRE�p��[�IF@Q���NACa%�$_}GœSTATUv�<œy�MAILAb�1x�!
�5�LAST�!��1"$ELEM_�� �\�iFEASIl3�nbg�Z�2�� >�96���`�pI�����G"�Q=� ��n2AB$U�0E���PV�!�6�BAS�2�5�r�AU8�P�PJ�$�1�7RM�@Rh3Ł���3`���P�r�!�4 ��$"S�~�	E2 2� �c���d +F�2*G�2"Э`���28VGW�DOU�����r�"$P �@�)G�RID��U�BAR�S�WTYm�"OT�O����� t�_"�$!��B�DO��\�� � ����P�OR���C���CSReV� )TVDIS�T_�P4PFT�PPW�P�PW4NY5NY6NY7�NY82Qn�Fbr_�~r�$VALU�3�(�+4j�A�F[��� !h^����C�!%���AN'��R�!���T")1TOTAL�_�$l06bPW=#I|�AKdREGENIj^b��X�8��=�� f� �TR�3�"Ia_S+��g^`��V���b��2E�# �?�(2��� cV_H�@DA8 ��`pS_YY����a&S8�AR �2�� �IG_SE�6�`R�%_���dC_�F$CMm�f�wrKDEh�?p�rI]��ZvsPsq!�F��H�ANC&�� p�Aj�"d#qIN�T1P��F}���M�ASK퓸0OVR ��� �<�!Ł�Gy��S�E�d�OJ6�k�F��PSLGHp�Q� \ 1�b%Z�$��3`� S���$�q�UY�y����c��ZQU�n�w�TE��@�' (�aJV�Q��q#IL_Mp$�Vt2����TQ ���R�0C���VB�CP��P_�J�Z�Mq�V�1p�V1~�2��2�~�3��3~�4��4 ~�� ��<�����;IN�VIB0�J��7��>�2:�2F�3*:�3F�4:�4F��� Y�r�U��gP
�tP���'��PL� TOR$��IN��u��5����T $�MC_FC�X�B�LC�B��u)`M��1I�s*�rC ��)���r��KEEP_H/NADD#�!e��0o�C�ѳ����A$�����O�d�>"��`����w��REM��@���!�Bµٱ޸U�$�e��HPWD  ;e�SBM�q�@?COLLAB"��Ph��'a�" IT' ��INO)�FCAqLh�
���� ,���FLnб1$SY�N���M��Ccr�~�`UP_DLY��=�r�DELA���!Z�"Y �AD �.��QSKIPG�� 	�
P��O��˂K���P_����Ƕ��� ��#ٖ#�gP"�tP "ځP"ڎP"ڛP"ڨPz"�9��J2R *���dX�0TJ#�� ��)1�Ѭa�����a�� RDCaw�� %�� R��R�!�8=��-DRGE� W3�{BFLG�0��sSW{	-DSPC���!UM_����2T�H2NuA��� 1�  ���|�A[ � D��x�x]�02_PC����S���1Q L10�_Co"/����q ���JPٰ7��6�K�+��� �.� NE���N���b\r�3�k����p����D�ESIG��JEVL�1��1��k��10Nٰ_DS�K�����EFC11��� �lV�������iI�AT����AS'J N�$	C�
���HGOME4����2������� 2D 
��3���gy����� ��4�����,>�5���as����
V6�����//(&/8/�7���[/m/0/�/�/�/ x��8����/�/�/? ?�2?PS)�����@�1��s`Y�V۰E�D� T���4,f�3�IO��
II�0XrOe�_OPE.C&b�3ަ�POWE��� �0����NK���&d �}�eB$wDSB��GNAr��%c��C��t��S2;32�5� ��Z5���׀ICEUS�/cSPE���QPA�RITq$aOPB�Q��RFLOWApT�R�01b�UJsCU8�@6��QUXT�q�Q>�pERFAC�Dʰ�U `VSCHN�Q� tV��_�@�kpc�$�`�`OM�*p��A>�#�p%�UcPD<����aPT�0F|uEXЙX|S!%��FA?��rj�r�a �� ���`;b K�AL$� ��U���]B�a  2� ��S���0�	Ч �${�����G+RO�`*dT�(p�6fDSPBfJOG@�`�C����AZ�N�������"VK�P_McIR^a~d�MT3��cAP%����`}t��Sp�`R��
��e�BRKHUQ�V��A;XI�1  �bc��r-b�q9�7e�`BS�OC6f۰N2uDU�MMY16O�$�SV��DE3A�CF��wK�0�D�pcOIR{ws0N�p|vFpl�w[`OV^eSF�z'RUN�s�rF�vQނcUFRA�zTO�TLCH�����OVlt[�[`WP�7�[c����r?p��_�p�� @h�TINVE\G@n1OFS\�C�P�WD�q��q>qf2,�eXpTRr��1a��E_FD�aMBS_CW���B��B�@*��ałˁ?�epV9Q ��P&��írGƇ�hAM�c��VP�F�!��_M݀R_�CS�T�$����Q�3T$HcBK�Q�fm�IO�5q|�&A��PPAp����������,�&BS�DVC_DBъ0ސ �Q�Bސ7�Q������F���3��L�E���+Pĉ`lqU�3P`FCAB�Ё2~㷀8û` �ڋ�O�UX�fSUBCP�[�-��/� �P/Ѯ�ރ�bB~��$HW_C�� 	P/ы��?�q0#�N�P�$UP�t	�>�ATTRIh���h`CYC��g�CA�B��cFLTR_2_FI�3�IH��F���PtkCHK�_S�CT�cF_�F_����FS�A��CHA�}�ֱ�RղRSD���Aq�S�A&@_T�}�.����PEM�0��MsT�ò/��Pò��K�D�IAG�URAIL�AC듑�M`LO�"p��Hv_�$PS�Nb�2 �L��PRRߐS}�I���Cё�f�	E�FUN��*QRIN1�}�|0^���Đq�S_;`���X����0f���P�f�C#BL���.�A'�#�*�#�DAp��h�.�'�LDyP`p����Ca2�����TI�°����P$CE_R�IAa�BAF��Pb�A��~���T2}�1C�S�؁OI���DF_L�0�r�Q�P�LM�F^�HRD�YO�af�RG��H����a|0p�/�MUL�SE�����Qp��$JxzJ�r�w�{F?AN_ALMp����WRN��HARDH�0�VZ0P]R�2����A��e_��fAU��RȴRTO_SBR&E�O`#��ӓ|��;�MPINFQ���N��Y�REGF�6NV�Pf3�fDA@�N��FL��R�$�M�Ѕ�`S����Pl����CMѐNF-�F�1����h��A��0;$�1$Y oQ�b�Q�0�� ��cEG�0+c`p�+AR=`CHu25pRr:T��eAXEEgwROBBjREDBf�WR,� q_�$sS�Y�`ep�S�WcRI,�>�STr@PCcPp�pE��0"G6Rr��;`B� R�r�7��2�OTOi�9�0��ARYBc40~�2��2t`FI�`�c�$LINK�GkTHS�PT_��R�F8Rr|XY�Z�R�9�OFF�Z�S{o8B@`���/��@�P�FI1�����CXt��Zd_J�A�R�r`0����30Rr�@��*!m�b"CFA�eD�Un�Hu3����TU�R��X�ӛ%BI�X� `�J'FL|�a�P8 � ��	3ʡg�� 1��0Kg`M �d�&Qs�����°�pSORQ&�Oa�P(���`O� �1ɐj4��Ma���~4OVE�1M IPk1��5�5�6�_Q�7c��7��4AN ڡV�1���1�`�0 �k1�5�1�7(E(EL�3OaERla�	��!E,��P��fDAA�P���!�@o�l�o�AX/��Ro�2��U �EQ��I{��I���JN  �J�J$�J��J��J1[ �F/��I/��I /��I/��I/�Y/�Y /�(Y/�8Y/�HYeQYYoDEBUڣ$��`��U�	ao�wABo��m��q3Vb�٢ 
$b�LeʡXgQq Xg��XgNXgXg$ Xg�Xg���g ��U.�LAB�J5֠��GRO[�J"��K�B_/�MF��s�� �v5qK51u�=vAND0��[DL��^A�zw K���� �x1��xN�NT��#��pVEL5��4�qm��xl9��NA��k ��$��ASS  �����* f*  �_�SI@���#���)�IY�n��(�AA{VM��K 2 T�� ?0  �5���r������ ��A	݀΍�* U��ߏ��!�͌@�L�܁`R�������e�BS�1�  16�� <u����
� �.�@�R�d�v����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶����� �����"�4�F�X�j� |ߎߠ߲���������ܱ��pMAX/� v���ʓ  d��IN�*��PRE/_EXE;�g�J��!43��T�e�IOC�NV�"<� �&�P���a ;�Ɨ��IO_�� 1r�P $�b�����V���U�?�����$�6�H�Z� l�~������������� �� 2DVhz �������
 .@Rdv�� �����//*/ </N/`/r/�/�/�/�/ �/�/�/??&?8?J? \?n?�?�?�?�?�?�? �?�?O"O4OFOXOjO |O�O�O�O�O�O�O�O __0_B_T_f_x_�_ �_�_�_�_�_�_oo ,o>oPoboto�o�o�o �o�o�o�o(: L^p����� �� ��$�6�H�Z� l�~�������Ə؏� ��� �2�D�V�h�z� ������ԟ�����LARMRECOV ~�!�J���LMDG ����� �LM_IF ��+��ߥ��� ɯۯ骓���0�B�~S�, 
 S� |��������ƿؿ�$�����1��U�g��yϋϝ��NGTO�L  ~� 	 A   ������PPINFO Z� Y��*�<�N�!�  f�P�~� ?�mߧߑ��ߵ����@��%��5�[����� ��������������)�;�M�_�m�PP�LICATION� ?����g�Han�dlingToo�l �� 
V9.10P/30���j�
88340̯���F0����10�28��������7�DF1��j���No�nej�FRA�j� 6w�_�ACTIVE� � ����  �U_TOMOD� ^���ÊCHGAPO�NL� �OUPLED 1��� 
 2��CUREQ 1	���  T<<�<	����@�w<���ƂHk�HTTHKY�A�o ���////�/S/ e/w/�/�/�/�/�/�/ �/??+?�?O?a?s? �?�?�?�?�?�?�?O O'O�OKO]OoO�O�O �O�O�O�O�O�O_#_ }_G_Y_k_�_�_�_�_ �_�_�_�_ooyoCo Uogo�o�o�o�o�o�o �o�o	u?Qc �������� ��q�;�M�_�}��� ������ˏݏ��� m�7�I�[�y������ ��ǟٟ����i�3� E�W�u�{�������ï կ����e�/�A�S�0q�w��NTO�����DO_CLEA�N���NM  �� <_�q���ϕϧ�BDSPDgRYRϊHI� ;�@L��%�7�I�[� m�ߑߣߵ��������MAX~�������	�X���PLUGG� ����PRC��B9�"=����c�Oh���^��SEGF� K�� ����9�K��%�7�I�8[�����LAP��� �����������	�-?Qcu��T�OTAL+�T��U�SENU��� �޸��NRGDI_SPMMC��0�C���@@���O�������_STRING 1
��
�M� S��

^_ITE;M1h  n�� ������// &/8/J/\/n/�/�/�/��/�/�/I/O SIGNALb�Tryout� ModeiI�np0Simul�atedmOu�t,<OVER�R�� = 100�lIn cyc�l 5mProg� Abor63m~4Statusk�	Heartbe�atgMH F�aul�7�3Aler�9�/�?�?�?O#O�5OGOYOkO}O  ��d��v�O�O�O�O __(_:_L_^_p_�_ �_�_�_�_�_�_ oo�OWOR��dJa�O $oro�o�o�o�o�o�o �o&8J\n������~PO b�1�pbk��#�5� G�Y�k�}�������ŏ ׏�����1�C�U�g��rDEV�~��� ���˟ݟ���%� 7�I�[�m���������ǯٯ����PALT�M6�bo�^�p� ��������ʿܿ� � �$�6�H�Z�l�~ϐ���$�GRI�d�� N�����&�8�J�\� n߀ߒߤ߶������߀���"�4�F���� R �M~���X������� �� ��$�6�H�Z�l� ~�������������l�PREG:�# ���� J\n����� ���"4FX�j|��-�$AR�G_J`D ?	�������  	$��&	[�]����')�SBN_CONFIG� �$1�#2=!!CII�_SAVE  ��$F!9#�TCEL�LSETUP ��%  OME�_IO�-�,%M�OV_H� �/�/R�EP���/�UTO/BACKv!�@"FRA:\� �/F '`r�0C8� T;�?  23�/07/18 17:50:04(�?�?�?�?4<��O6OHOZOlO~O�O�$O�O�O�O�O __�O<_N_`_r_�_ �_�_3_�_�_�_oo &o�_Jo\ono�o�o�o\�o���  /1_3�_\ATBCKCTL.TM���op+=;INI9��v56%J!0MESSAGV dqF!�o{ODE_D� Y&6%��xO���3PA�US� !�� , 	� x���,		� 8�"�\�F�X���|��� ���֏����F���t�pTSK  ��}C?I0UPDT̝pbwd���vXW?ZD_ENBbt2*��STAau�����XIS$ UNT �2�C!E � �	 8�� �����!D �� �p� �/Q"
���.������
9�r����F�Е��/6�5��5 [?^. 8��a�¯p��������MET��2i�b# P�B���A�-mA��J 7MWAA%��A��٭�>a:>ٻ��>p�35ؔ�>B�>H�0��SCRDCFG� 1�%1 �^%C"篻�Ϳ@߿���<?
QZ) ��e�wωϛϭϿ�&� ��J���+�=�O�a�0��߼1GR���X����`NA� �s	4��_ED`p�1���_��%=-�`EDT-���*H�B�Y�b?$� -3�
"O�&
�^��  ����2��#� �G��_���G� ���6����3��+ ]���̔\��Z�l�����4K����� ��t�&8�\��5�d���@� ��(��6�S 0/w��/w/��f/���7�//�/C/����/C?�/�/2?�/��8{?���?�f&��?O V?h?�?�?��9GO�?�O�?i&�pO�O"O4O�OXO��CR���/__ q_ =:_�_�O�O�_"_�����NO_DEL��ߞ�GE_UNU�SE�ߜ�IGAL�LOW 1���   (*S�YSTEM*֣�	$SERV_GqR�k_`�pREGhe�$�c֬_`NUMx�j�c�mPMU`>֥LAY�֬�PMPAL<ap�eCYC1p��c� }�`�n%sULS�U�o�mr�qjcL�;ttBOXORI��eCUR_ap�m�PMCNV�f�ap10~�pT4D�LIǐZ|i	*P�ROGRAgdPG_MI�n�)��AL�u6� �)�B�T�_n$FLUI_RESUw���o���ÄMRvn�`�\ �_Β��+�=�O�a� s���������͟ߟ� ��'�9�K�]�o��� ������ɯۯ�����#��RLAL_OU�T Nk���W?D_ABORp/o���ITR_RTN�  �D��ل�N�ONSTO�Я�� 8hCE_RIA3_I,`��������FCFG ����ĨN�_LI�Mvb2�� �?  � 	��gϢ�B<�҄��e�@�� VϷ����ϨH
���ߒ�2�PAn�G�P 1��ޥ�n߀ߒ�Q�C>�  C.���f��z����߶Ї�Б�Ж*�Р�Ъ�д�Թ�`����������C���_ǀ CѶ��J�m�G?��HE�P�ONFIπ��d�G�_P�p1;� �U;ծ������������,�d�KPAU�S~q1;���  �r.�t�;�b������� ��������0@�fL����6�M~��NFO 1?�;� �T���B�̵���5Au�9	��]�Ǝ�@���K D5O�y���C����($6�T�5+��P�� 8�h�Ca���.~:���1５��O��ϨG��CO�LLECT_�0?�x�ǯEN�p�������NDE��?�;c�R12�34567890�'�Bya�//&��HC��C)j/�/y\i/{/ �/z[�/�/?�/�/? `?+?=?O?�?s?�?�? �?�?�?�?8OOO'O �OKO]OoO�O�O�O�O�_�O�9�� ���IO !)������_�_�_l�_`WTR6�2"D]�(�{Y
�O�^o��#o] jt�i_MO�R9�$;� ��:B��\`�e �i �o�o�o�o�o�kbb1�*:�%pm,t�?]�]�H��>q�KFt�`�R�&�utqtrC_4  A�����Mx�A����B�p�Cd B��d C � @�r��q�:Sd�QbZqI#'d}�?�s9�(pm����d�ZqT_DEFB� �{%oR��thPN�USE��s���g�K�EY_TBL  �������	
��� !"#$�%&'()*+,�-./(':;<=�>?@ABC)�G�HIJKLMNO�PQRSTUVW�XYZ[\]^_�`abcdefg�hijklmno�pqrstuvw�xyz{|}~����������������������������������������������������������������������������,���͓���������������������������������耇����������������������4Q��LC�Kp�ٹ��p�STA����t_AUTO_�DOζkv�IN�D�ٞ�R_T1���T23�ݵʳ���TRL(�LET�E��z�_SCR�EEN ;�_kcsc�Uʰ�MMENU 1)l� <7�@���� ��F��#�I���Y� k��������ſ׿�� 6���l�C�UϢ�y� �ϱ������� ���	� V�-�?�eߞ�u߇��� �߽�
������R�)� ;��_�q������ �����<��%�r�I� [��������������� &��5nEW� {�����"� X/A�ew�����/)\ʠ_M�ANUALo�*�D�B'a.b����DBG�_ERRL.�*֫�Q /�/�/��.L!NUMLI�M���lu
L!P�XWORK 1+֫�/#?5?G?Y?k?�mDBTB_�� �,{-�s�Qst�3QDB_AWAYzT#�QGCP lr�=���"�2_AL� ٟ�2P"Yn���lp�E(_n  1-�[,p
?POJf@O}O�6�_M�IS֐�;@|�p�CONTIM����lt��FI
�� CMOTNEN�Dt�DRECOR�D 13֫ �<�OxsG�O�KQ9_ x{�2w_�_�_�_DX�_ �_K_ oo_$o6oHo�_ �_~o�_�oo�o�o�o �o�o �oD�ohz ���1�U
� �.�@��d����� ����Џ�Q��u�� ��N�`�r���󏨟� ��;����&���J� 5�C������ȯ7� �ׯm�"���F�X�j� �y����Ŀ3���� ϣ���Bϱ�f�տ�� �Ϯ���[���S��w��,�>�P�b��Ͽ2TO�LERENC�4B��B�0L��L C�SS_CNSTC�Y 249�Y e�B���������� #�5�G�]�k�}��� ���������������DEVICE 25�� �6o��� �������������&�O��HNDGDg 6�۬0Cz9
|Q��LS 27Y�8������:��PARAM 8,I�2�5&��ySLAVE �9YE_CFG �:F&dM�C:\��L%04�d.CSV%@c��B�A �CH kkO&/B/X�&2"_!o/])\!1@JPя#N.A��1n_CRC_?OUT ;Y��1~*_NOCODz�<,G�SGN �="UR#M��20-JUL�-23 02:5y7�0A18>5�17:51�~�? V�hr9n1�&o061�M��?Þ�j��1�>��VERSION� ):V4�.2.11�KEF�LOGIC 1>^�� 	�(1@�I�!M�2PROG�_ENB Xa=CU�LS�G `�2_�ACCLIM�F����|CWRSTJNT�G
S�ц�1MOFLX!2�DI?NIT ?��"Uv�� �FOPTu� ?	�F�B
 ?	R575&'P�74,Y6-X7-W50QX�4WR2-T�({_|�7
TTO  ]�?�_�6V�@DEXҩGd�B� �SPA�TH A):A�\�_5oGo|�HCP�_CLNTID y?�6� �+�Ӈo��IAG_G�RP 2D� �� 	 �D�  D�� �D  B��Т��ff�j�`���oĝl�a���%���B�N�C�-Bz��Bp���e`�imp�2m7 7890?123456xq�G��`�  Ao��
Aj{Ad��]AW��AP��AJ=q�AC33A<�4cz�j�p�!@���]pA�q��A��,���B4�lf�d�X�!
�ru�ppQ��Aj�HAeG��A_�pY��A�S�pM2�F�RA@(��J���t�Jx��I�@�p���������@��H�L�^�p��������3�3<��=q@~��R@xQ�@q���@k�@dzw�@]��Vff؏����� ���s>�l���@e@^�J�W
=@Pv�G��@@v�7ڐ.{d�v����������S>�M���AR�<�(�@5Ґ/\)�@(��@!R� ֏ ��$�6��ĭ� ��ܯ"�4����V�|� Z�����<�N������ �0�B�̿R��B�`�r�5���M�ّe��m>���R��?�33?�9������m7'�Ŭ��6��4�F���L�m@�T�����ڐ␀N��Њ=@�pAh������c= c<���]>*�H>�V>�3�>�����m<����<b�a�i�L. ��?� �C� � <(�UX" 4�>��ё��ٝi	A吳 ?�el���t� ���,��H��8�b����r��z����x�?��7��>�(�>�!����=�����m��G��G�@�m����I��m�����i�@�Ҁ�@Q�?L��Ly�o�g�v(\����]p'�@�����8���	�gC�> ���Cu��<Zl <� ����`��&%��18� �����4J6�<��D5OL��rC��� �5�q�W�S����$�z�	�($6�T��Á� i��x��������ʝm;���t��9/�aCT_�CONFIG �E?i3eg��%�aSTBF_TTS�G
UI�#�0�Ct�A�&� MAU�@�JOJ"MSW_CF�X F�k  �p�:O�CVIEW� G�-�a���o=?O?a? s?�?�?�B+?�?�?�? �?OO�?>OPObOtO �O�O'O�O�O�O�O_ _(_�OL_^_p_�_�_ �_5_�_�_�_ oo$o �_HoZolo~o�o�o�o Co�o�o�o 2�o�Vhz���@,RC�#{��"!L�~� ��A�0�e�T����$�SBL_FAUL�T I�z 8��G�PMSK�'��L TDIAG J\)��!��1��UD1: 6789012345�p"1�j'�uP&/O�a� s���������͟ߟ� ��'�9�K�]�o������y��
>���F&TORECP���
� ��%���=�:�L�^�p� ��������ʿܿ� � �$�6�H�Zρ��������7UMP_OP�TION� ����T�R�"�#����PM�E�%��Y_TEM�P  È�33BȞ 1��A.�ԇUNI� �%1��&Y�N_BRK K�?6EDITOR�����
��_ԠEN�T 1L�y � ,&PART1 TLOG �����f���2���&�MAI���߫�?&OMAY��[� ��F��߇���� u����J�����
IRV�WAI����&-�BCKEDT- ���/���PICKSIM_��[���y���o"�x������� ������3Wi P�t�������~�MGDI_�STAD� !1�y�N�C71M�+ �P`�r��
��d�� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?��j? |?�?�?�9��?�?�? �?
OO.O@OROdOvO �O�O�O�O�O�O�O_ _*_<_�:c?m__�_ �_�?�_�_�_�_o!o 3oEoWoio{o�o�o�o �o�o�o�o/A [_ew���_�� ����+�=�O�a� s���������͏ߏ� ��'�9�SA�o��� �����ɟ۟���� #�5�G�Y�k�}����� ��ůׯ�����1� K�]�g�y���A����� ӿ���	��-�?�Q� c�uχϙϫϽ����� ����)�C�U�_�q� �ߕ߯���������� �%�7�I�[�m��� ������������!� 3�M�W�i�{����߱� ��������/A Sew����� ��+E�Oa s�������� //'/9/K/]/o/�/ �/�/�/�/�/�/�/? #?=/?Y?k?}?�� �?�?�?�?�?OO1O COUOgOyO�O�O�O�O �O�O�O	__5?G?Q_ c_u_�_�?�_�_�_�_ �_oo)o;oMo_oqo �o�o�o�o�o�o�o �_?_I[m�_ �������!� 3�E�W�i�{������� ÏՏ�����7A� S�e�w��������џ �����+�=�O�a� s���������ͯ߯� ��/��K�]�o��� �����ɿۿ���� #�5�G�Y�k�}Ϗϡ� �����������'�9� C�U�g�ߓ��߯��� ������	��-�?�Q� c�u��������� ����1�;�M�_�q� �ߕ����������� %7I[m� ������)� 3EWi����� ����////A/ S/e/w/�/�/�/�/�/ �/�/?!+?=?O?a? {m?�?�?�?�?�?�? OO'O9OKO]OoO�O �O�O�O�O�O�O�O? _5_G_Y_s?�?�_�_ �_�_�_�_�_oo1o CoUogoyo�o�o�o�o �o�o�o_#_-?Q c}_������ ���)�;�M�_�q� ��������ˏݏ�i %�7�I�[�u��� ����ǟٟ����!� 3�E�W�i�{������� ïկ�����/�A� S�m�w���������ѿ �����+�=�O�a� sυϗϩϻ������� ���'�9�K�e�[߁� �ߥ߷���������� #�5�G�Y�k�}��� �����������1� C���o�y��������� ������	-?Q cu������ ���);Mg�q �������/ /%/7/I/[/m//�/ �/�/�/�/�/?!? 3?E?_i?{?�?�?�? �?�?�?�?OO/OAO SOeOwO�O�O�O�O�O �O�/__+_=_W?I_ s_�_�_�_�_�_�_�_ oo'o9oKo]ooo�o �o�o�o�o�o�O�o #5O_a_k}�� �������1� C�U�g�y��������� ӏ�o�o	��-�?�Y c�u���������ϟ� ���)�;�M�_�q� ��������˯E���� �%�7�Q�[�m���� ����ǿٿ����!� 3�E�W�i�{ύϟϱ� ���������/�I� S�e�w߉ߛ߭߿��� ������+�=�O�a� s����������� ��'�A�7�]�o��� �������������� #5GYk}������� �$EN�ETMODE 1�NB�� W �������� RROR_PROG %�
�%��an<TAB_LE  �L�����<SEV�_NUM 
  � <�_AUTO_EN�B  (9_;NO! O�} "  *�Y ��Y �Y �Y  +�X r/�/�/2$FLT9R/0&HIS����++_ALM 1]P� ���Y,��+�/2?D?V?h?�z?�?�/_�8   ��W!�:� T�CP_VER �!�
!Y�?$EX�TLOG_REQ��&�))#CSIZ\,ODSTKIIG%�� BTOL  ���Dz�"�A= D_BWD�0�@��&�A#�CDI�A ;QB��C<��KSTEP�O�O|� �@OP_DOkO��FACTORY�_TUN�'d3YD�R_GRP 1R�	�!d 	�?�_�{P�*u����RHB ���2 ��� �e9 ����V{S�_��]{PB���B��F>C��B����AԂ=Bu�� �[A���B��B��A����AI��B ��]�_WoBo{o�fo�o�o�o�o  @��:A|=@�9q��o��
 �F�5W&b�`��A�$� #�4<�o`�K��Y�  �qAݠ�`�33�r�3�3�]@UUT�z@��`�pj$>u.��>*��<�����]E�� F@� �p&��]J���NJk�I'P�KHu��IP��sF!���]?��  j��9�<�9�89�6C'6<,�5���~����=����a��� �_&����#tFEATU�RE SB��@�"Hand�lingTool� 	���Eng�lish Dictionary��4D St��ar�d	��Analo�g I/O@�I�g�le Shift�\�uto Sof�tware Up�date��mat�ic Backu�p���groun?d Edit���CameraW�F�[�CnrRndI�m���ommon� calib U�I��n͑�Mo�nitor&�tr~�Reliabp���DHCP�]�a�ta Acqui�s5�^�iagno�s��T�x�ocum�ent View�eA�`�ual C�heck Saf�ety!��hanGced!����sʠ�Frސ�xt. oDIO 1�fi���&�end��Err�@�L��B��sA�r�R�1� �@�FCT�N Menu�v|\���TP In���fac���Gig�E��εƐp Ma�sk Exc��g�#�HT��Prox�y Svˤ�ig�h-Spe��Sk�i�Ŧ�5�mmuwnic��ons<ȃur����s�X���c�onnect 2�s�ncr��str�u#�qʚ�e��۠J����KAREL �Cmd. L �u�a���Run-T�i"�Env�Ȅ�e�l +��s��S/�W�Licens�eݣʬX�Book�(System)��MACROs,~3�/Offsew��V�H5���q�[�MR�:�6���MechStop�t����V�iS�s���x��T������odq�witc�h�ߚӡ�.{��O�ptm,���fi�lʬ��gi�V�ul�ti-T��Г�P?CM fun�Ǣ��o��ޢ����RegeiK�rW���rià�F����U�Num �Sel��� � AdjuG��=�s�N�tatu��f�Ū��RDM Robo}t �scove)���ea��"�Fre�q AnlyW�Rem��5�n7�����Servo5���?SNPX b�x�;SN��Cli¡%t�Libr(�E��Q ��W o0�t���ssag����0 0��n���0/I����MILIB��P� Firm���PΡ�AccǐϛTPsTXm��elnn�����jղorq}uq�imula?�4�bu�Paѱ�ƐZ�(�&�ev.̞��ri۠:U�SB port ��iPL�aà�R� EVNT��n?except���������VC�rR�I���V��o"�%4Wz+S8 SC4�/gSGE�/�%UI�?Web Pl}� >�i�'4�����x�ZDT ApplP���&?|7Grid��playv=� ��
�7Rf".7��6���/�Y�-10iA/8�L�?Alarm Cause/���ed*�Ascii<�<�Loadʠ:J'UplP@�l�7�#Gu=�rO�BP��Ֆycp�����蠕��RA� �9�NR�TJ�On�e Hel��漿�������1tr;�ROS� Eth
�t�Be�W7iR�$2D PYk;�uVIm+�Fd�� �^nsp���Q��64MB DRA9M�O�SFRO�_ېgellW��shaDo gcK�e��p�2ltyp�s'�ԗ�Bt��D�.�maiܠ�;�T�qV�Rt7��FL!PSup��c��� pL���cro�~���W�4��&��au7estz&rtڡ���/�3DL}|�Q����Ty,K��l B�ui��n�/APL�C��uVZ��/CG�l��CRG#��$D���@�R�LS[��%B�Uw��%Kі��!T	A���B�,يE�TCB��ʏ��/��^�TC��v�8�%��TEHǟٖ�"�ؗV�����/��F�H����G:���n�Ȁ�����H¯��IA0߯�ޯ��LN����M��D���D�����N����P��������R�R���Sڿ�����Wp.�@Ǣ��$VGFf�x�P2Z���2��ǂϒ��B�ϔ�D�ϔ�Fpr�����"TUT�01J�\�2f�\�T�BGG��rai�n��UI*ЦUHM9I��r ponU2�8����af{ �R�v�VK�AREL��_TP� �e��R9�0�B� o�f�x�������� �����5�,�>�k�b� t��������������� 1(:g^p� ������ - $6cZl��� �����)/ /2/ _/V/h/�/�/�/�/�/ �/�/�/%??.?[?R? d?�?�?�?�?�?�?�? �?!OO*OWONO`O�O �O�O�O�O�O�O�O_ _&_S_J_\_�_�_�_ �_�_�_�_�_oo"o OoFoXo�o|o�o�o�o �o�o�oKB T�x����� ����G�>�P�}� t�������׏Ώ��� ��C�:�L�y�p��� ����ӟʟܟ	� �� ?�6�H�u�l�~����� ϯƯد����;�2� D�q�h�z�����˿¿ Կ���
�7�.�@�m� d�vψϚ��Ͼ����� ���3�*�<�i�`�r� �ߖ��ߺ�������� /�&�8�e�\�n��� �����������+�"� 4�a�X�j�|������� ��������'0] Tfx����� ��#,YPb t������� //(/U/L/^/p/�/ �/�/�/�/�/�/?? $?Q?H?Z?l?~?�?�? �?�?�?�?OO OMO DOVOhOzO�O�O�O�O �O�O_
__I_@_R_ d_v_�_�_�_�_�_�_ oooEo<oNo`oro �o�o�o�o�o�o A8J\n�� �������=� 4�F�X�j�������͏ ď֏����9�0�B� T�f�������ɟ��ҟ �����5�,�>�P�b� ������ů��ί��� �1�(�:�L�^����� ������ʿ��� �-� $�6�H�Zχ�~ϐϽ� ����������)� �2� D�V߃�zߌ߹߰��� ������%��.�@�R� �v��������� ��!��*�<�N�{�r� �������������� &8Jwn������  ?H552���21R785�0J614AwTUP)545)�6VCAMC�RIdUIF)2�8eNRE52�XR63SCH�DOCV�CS]U869)04�EIOC�4R{69XESETAvWJ7WR68�MASKPRXuY}7OCO(�3A! (3`&J�6'53�H�(L{CHH&OPLGA�0x&MHCRI&S��'MCS@0$'5=54MDSW!7k';OPk'MPRl&���(0(PCM|R�0g7! 4� �'51�L51�80LPR�S'69`&FRD�dFREQMC�N93(SNByA��'SHLBF�M'G�82(HT=C@TMIL��TPA�TPTXFYFEL�6� �8�J95�TU�Tl'95`&UEV�&UECH&UFR�dVCC XO�&V�IPdFCSC�FC�SG��IWE�B@HTT@R6l��HCG_WIGGWoIPGS�VRCdF�DGk'H7�R6�6LR7'R�8R[53�768�82x&�R�*4�W664R�64NVD&R�6�'9 �X�9 �Du0+gF~hCLIP8�KCMS��`@S�TY$WTO@NN�`&ORS�&M�8O]L�hENDLW�S�hFVR�V3�D$X{PBV�FA�PL�APVl&C�CG@CCR�&C�DWCDL�VCS�B�CSK,6CT�{GCTBHV�p�hCh(F�p�xC<WTC|l�ppwTC�wTC&�CTE�9�|wTEX�9�0WTF�xF�h�G�xGx�$�H$�IpF��$��GCTM�hUM�M�xN$�P��eP�xR�x�hTS�x�W8��VVGFP�P�2 WP2�6e�\�Bj\�D\�F|VP���VT��VTBZ�wV�IHWGV�P
՗K$WV_V��)� ;�M�_�q��������� ˯ݯ���%�7�I� [�m��������ǿٿ ����!�3�E�W�i� {ύϟϱ��������� ��/�A�S�e�w߉� �߭߿��������� +�=�O�a�s���� ����������'�9� K�]�o����������� ������#5GY k}������ �1CUgy �������	/ /-/?/Q/c/u/�/�/ �/�/�/�/�/??)? ;?M?_?q?�?�?�?�? �?�?�?OO%O7OIO [OmOO�O�O�O�O�O �O�O_!_3_E_W_i_ {_�_�_�_�_�_�_�_ oo/oAoSoeowo�o �o�o�o�o�o�o +=Oas��� ������'�9� K�]�o���������ɏ�ۏ�  H55Ȕ������R78�50	�Jw614	�ATU��?�5459�6	�VwCAM	�CRI���UIF9�28��N�RE�52x�R6�3�SCH	�DO�CV��CSU�8�699�0H�EIOuCɛ4(�R69x��ESETY�w�J7�w�R68�MAS�K	�PRXY��7.	�OCOy�3Y�(����8�3تJ67�5u3(�H�LCH���OPLGY�0��M�HCR��Sw�MC�SX�0��55H�MgDSWٻ�OP�GMPR��(�08�7PCM��R07˅��H���(�51h�51�x�0h�PRSx�6�9تFRD��FR�EQ�MCN	�9=38�SNBAٛ�/SHLB	�M7�吺ȼ28�HTCX�T�MIL�(�TPA�H�TPTXy�EL��ʅ�(�8'�%��J�95��TUT�9�5تUEVx�UE�C��UFR��VCuCX�O��VIP��wCSC��CSGȚ��I	�WEBX�H�TTX�R6ל��C�G��IG��IPGmS	�RC��DG竻H7'�R66h�Ru7g�Rv�R53h˫68h�2��R6�4v��66H�R64�7NVDx�R6�����h�������D0��F�VCLI�g�CMqSH�� X�STY���TOX�NNتOR�S��M��OL�E�ND�Lg�S�F;VRH�V3D�짛wPBV��APLH�wAPV�CCGX��CCRx�CDg�C�DL(�CSB�C�SK�CT��CTB�� �C8�5 ,�C��TC��5 �T�C�TCx�CTE��� �TE�� ��TF,F�G,G�-�,H�,I�E0�,���CTM�Mx,M��N�,PH<P,R,,�TS,W�=(��VGFKP2X�PQ2��5@(LB(LD(LmF��VPW;VT�\�@(�VTB�V�KIHw�V5��KK��V���_1_C_U_g_ y_�_�_�_�_�_�_�_ 	oo-o?oQocouo�o �o�o�o�o�o�o );M_q��� ������%�7� I�[�m��������Ǐ ُ����!�3�E�W� i�{�������ß՟� ����/�A�S�e�w� ��������ѯ���� �+�=�O�a�s����� ����Ϳ߿���'� 9�K�]�oρϓϥϷ� ���������#�5�G� Y�k�}ߏߡ߳����� ������1�C�U�g� y������������ 	��-�?�Q�c�u��� ������������ );M_q��� ����%7 I[m���� ���/!/3/E/W/ i/{/�/�/�/�/�/�/ �/??/?A?S?e?w? �?�?�?�?�?�?�?O O+O=OOOaOsO�O�O �O�O�O�O�O__'_ 9_K_]_o_�_�_�_�_ �_�_�_�_o#o5oGo Yoko}o�o�o�o�o�o �o�o1CUg y������� 	��-�?�Q�c�u����������Ϗ���STD�LANG�� �2�D� V�h�z�������ԟ ���
��.�@�R�d� v���������Я��� ��*�<�N�`�r��� ������̿޿��� &�8�J�\�nπϒϤ� �����������"�4߀F�X�j�|ߎߠ߲�R{BT�OPTN�� �������#�5�G�Y�k�DPN����� ����������%�7� I�[�m���������� ������!3EW i{������ �/ASew �������* �/1/C/U/g/y/�/ �/�/�/�/�/�/	?? -???Q?c?u?�?�?�? �?�?�?�?OO)O;O MO_OqO�O�O�O�O�O �O�O__%_7_I_[_ m__�_�_�_�_�_�_ �_o!o3oEoWoio{o �o�o�o�o�o�o�o /ASew�� �������+� =�O�a�s��������� ͏ߏ���'�9�K� ]�o���������ɟ۟ ����#�5�G�Y�k� }�������ůׯ��� ��1�C�U�g�y��� ������ӿ���	�� -�?�Q�c�uχϙϫ� ����������)�;� M�_�q߃ߕߧ߹��� ������%�7�I�[� m����������� ���!�3�E�W�i�{� �������������� /ASe�h�������99���$FEAT_�ADD ?	����  	�%7I[ m������ �/!/3/E/W/i/{/ �/�/�/�/�/�/�/? ?/?A?S?e?w?�?�? �?�?�?�?�?OO+O =OOOaOsO�O�O�O�O �O�O�O__'_9_K_ ]_o_�_�_�_�_�_�_ �_�_o#o5oGoYoko }o�o�o�o�o�o�o�o 1CUgy� ������	�� -�?�Q�c�u������� ��Ϗ����)�;� M�_�q���������˟ ݟ���%�7�I�[� m��������ǯٯ� ���!�3�E�W�i�{� ������ÿտ���� �/�A�S�e�wωϛπ�Ͽ��������D�EMO S   �N�D� V߃�zߌ߹߰����� ������I�@�R�� v����������� ��E�<�N�{�r��� ������������
 A8Jwn��� ����=4 Fsj|���� ��//9/0/B/o/ f/x/�/�/�/�/�/�/ �/?5?,?>?k?b?t? �?�?�?�?�?�?�?O 1O(O:OgO^OpO�O�O �O�O�O�O�O _-_$_ 6_c_Z_l_�_�_�_�_ �_�_�_�_)o o2o_o Voho�o�o�o�o�o�o �o�o%.[Rd �������� !��*�W�N�`����� ��Ï��̏����� &�S�J�\��������� ��ȟ����"�O� F�X���|�������į ޯ����K�B�T� ��x���������ڿ� ���G�>�P�}�t� �ϳϪϼ������� �C�:�L�y�p߂߯� �߸�����	� ��?� 6�H�u�l�~���� ��������;�2�D� q�h�z����������� ��
7.@md v������� 3*<i`r� ������/// &/8/e/\/n/�/�/�/ �/�/�/�/�/+?"?4? a?X?j?�?�?�?�?�? �?�?�?'OO0O]OTO fO�O�O�O�O�O�O�O �O#__,_Y_P_b_�_ �_�_�_�_�_�_�_o o(oUoLo^o�o�o�o �o�o�o�o�o$ QHZ�~��� ����� �M�D� V���z�������ݏԏ ��
��I�@�R�� v�������ٟП�� ��E�<�N�{�r��� ����կ̯ޯ��� A�8�J�w�n������� ѿȿڿ����=�4� F�s�j�|ϖϠ����� ������9�0�B�o� f�xߒߜ��������� ���5�,�>�k�b�t� ������������� 1�(�:�g�^�p����� ���������� -$ 6cZl���� ����) 2_ Vh������ ��%//./[/R/d/ ~/�/�/�/�/�/�/�/ !??*?W?N?`?z?�? �?�?�?�?�?�?OO &OSOJO\OvO�O�O�O �O�O�O�O__"_O_ F_X_r_|_�_�_�_�_ �_�_oooKoBoTo noxo�o�o�o�o�o�o G>Pjt �������� �C�:�L�f�p����� ��ӏʏ܏	� ��?� 6�H�b�l�������ϟ Ɵ؟����;�2�D� ^�h�������˯¯ԯ ���
�7�.�@�Z�d� ������ǿ��п���� �3�*�<�V�`ύτ� ���Ϻ��������/� &�8�R�\߉߀ߒ߿� ����������+�"�4� N�X��|������ ������'��0�J�T� ��x������������� ��#,FP}t ������� (BLyp�� �����//$/ >/H/u/l/~/�/�/�/ �/�/�/?? ?:?D? q?h?z?�?�?�?�?�? �?O
OO6O@OmOdO vO�O�O�O�O�O�O_|_2]  )X H_Z_l_~_�_�_�_�_ �_�_�_o o2oDoVo hozo�o�o�o�o�o�o �o
.@Rdv �������� �*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n��������� ȟڟ����"�4�F� X�j�|�������į֯ �����0�B�T�f� x���������ҿ��� ��,�>�P�b�tφ� �Ϫϼ��������� (�:�L�^�p߂ߔߦ� �������� ��$�6� H�Z�l�~������ ������� �2�D�V� h�z������������� ��
.@Rdv ������� *<N`r�� �����//&/ 8/J/\/n/�/�/�/�/ �/�/�/�/?"?4?F? X?j?|?�?�?�?�?�? �?�?OO0OBOTOfO xO�O�O�O�O�O�O�O __,_>_P_b_t_�_ �_�_�_�_�_�_oo (o:oLo^opo�o�o�o �o�o�o�o $6 HZl~���� ���� �2�D�V� h�z�������ԏ� ��
��.�@�R�d�v� ��������П���� �*�<�N�`�r����� ����̯ޯ���&� 8�J�\�n��������� ȿڿ����"�4�F� X�j�|ώϠϲ������������0�  1�6�L�^�p߂� �ߦ߸������� �� $�6�H�Z�l�~��� ����������� �2� D�V�h�z��������� ������
.@R dv������ �*<N`r �������/ /&/8/J/\/n/�/�/ �/�/�/�/�/�/?"? 4?F?X?j?|?�?�?�? �?�?�?�?OO0OBO TOfOxO�O�O�O�O�O �O�O__,_>_P_b_ t_�_�_�_�_�_�_�_ oo(o:oLo^opo�o �o�o�o�o�o�o  $6HZl~�� ������ �2� D�V�h�z������� ԏ���
��.�@�R� d�v���������П� ����*�<�N�`�r� ��������̯ޯ�� �&�8�J�\�n����� ����ȿڿ����"� 4�F�X�j�|ώϠϲ� ����������0�B� T�f�xߊߜ߮����� ������,�>�P�b� t����������� ��(�:�L�^�p��� ������������  $6HZl~�� ����� 2 DVhz���� ���
//./@/R/ d/v/�/�/�/�/�/�/ �/??*?<?N?`?r? �?�?�?�?�?�?�?O O&O8OJO\OnO�O�O �O�O�O�O�O�O_"_ 4_F_X_j_|_�_�_�_ �_�_�_�_oo0oBo Tofoxo�o�o�o�o�o �o�o,>Pb t������� ��(�:�L�^�p��� ������ʏ܏� �� $�6�H�Z�l�~����� ��Ɵ؟���� �2� D�V�h�z�������¯ ԯ���
��.�@�R� d�v���������п� ����*�<�N�`�r� �ϖϨϺ��������(�&�5�:�-�P� b�t߆ߘߪ߼����� ����(�:�L�^�p� ����������� � �$�6�H�Z�l�~��� ������������  2DVhz��� ����
.@ Rdv����� ��//*/</N/`/ r/�/�/�/�/�/�/�/ ??&?8?J?\?n?�? �?�?�?�?�?�?�?O "O4OFOXOjO|O�O�O �O�O�O�O�O__0_ B_T_f_x_�_�_�_�_ �_�_�_oo,o>oPo boto�o�o�o�o�o�o �o(:L^p ������� � �$�6�H�Z�l�~��� ����Ə؏���� � 2�D�V�h�z������� ԟ���
��.�@� R�d�v���������Я �����*�<�N�`� r���������̿޿� ��&�8�J�\�nπ� �Ϥ϶���������� "�4�F�X�j�|ߎߠ� ������������0� B�T�f�x������ ��������,�>�P� b�t������������� ��(:L^p �������  $6HZl~� ������/ / 2/D/V/h/z/�/�/�/ �/�/�/�/
??.?@? R?d?v?�?�?�?�?�? �?�?OO*O<ONO`O rO�O�O�O�O�O�O�O�__&_8Y�$FE�AT_DEMOIoN  =T�hP��=PPTINDE�X][lQ�PPIL�ECOMP T�����Q�kRKU�PSETUPo2 U�U�R?�  N �Q�S�_AP2BCK �1V�Y  �)9Xok%�_:o=P�P(oeo;U�_�o o �oDo�o�ozo�o3 E�oi�o��.� R�����A�� N�w����*���я`� �����+���O�ޏs� �����8�͟\�ڟ� ��'���K�]�쟁�� ����F�ۯj������ 5�įY��f������ B�׿�x�Ϝ�1�C� ҿg����ϝ�,���P� ��t���ߪ�?���c� u�ߙ�(߽���^��� ���)��M���q� � ~��6���Z������ %���I�[������� ��D���h�����
3t�Y�PP�_ 2�P*.VR:���*��������n PC���F'R6:�4�X�T|P|�y��_PI���*.F�q/��	�<,8�`/�STMk/�/"�/�-O/�/�H�/?�'?�/�/i?�GIFs?�?�%�?pF?X?�?�JPG�?�!O�%O�?�?qO�
JS{O�O��7C�OOO�%
JavaSc�ript�O�?CS��O(_�&_�O %�Cascadin�g Style ?SheetsT_���
ARGNAME�.DT�_��� \@�_U_�A�T�_�_�P�DISP*�_����To�_�QNa\oo
�TPEINS.X3ML�o�_:\�o]o��QCustom Toolbar�o�iPASSWOR�DSo��FRS:�\#�oD`Pass�word Configd���<� ���+�=��a� �����&���J�ߏn� �����9�ȏ2�o��� ��"���ɟX��|�� #���G�֟k������ 0�ůT���������� C�U��y������>� ӿb�������-ϼ�Q� �Jχ�ϫ�:����� p�ߔ�)�;���_��� ���$߹�H���l��� ��7���[�m��ߑ�  ����V���z���� ��E���i���b���.� ��R���������A S��w�*<� `���+�O� s��8��n /�'/��]/��/ /z/�/F/�/j/�/? �/5?�/Y?k?�/�?? �?B?T?�?x?O�?O CO�?gO�?�O�O,O�O PO�O�O�O_�O?_�O �Ou__�_(_�_�_^_ �_�_o)o�_Mo�_qo �oo�o6o�oZolo �o%�o[�o ��D�h��� 3��W�������� @����v����/�A� Џe�􏉟��*���N���r�������$F�ILE_DGBCK 1V������ �< �)
SUMMARY.DG#��ϜMD:W����ېDiag S?ummary�����
CONSLOG���p���ۯ���C�onsole l�og���	TPA'CCN�v�%^������TP Acc?ountin=����FR6:IPKDMP.ZIPϿ�Ә
� ϧ���Exception$��ջ��MEMCHECCK��������/��Memory D�ata����l{�)��RIPE�p�ϒ�'߶�%��� Packet yL<���L�$�e���STAT!��߾�� %C�S�tatus��`�	FTP�������1�mment �TBD4�`� >I�)ETHERN�Ey��f�w�瑱?EthernL�3�?figuraCϫ�~�DCSVRF(��� �9����� v�erify alyl<���M.c��DIFF1��)���<=�S�diff��t�|f���CHG01�������C����kv�- 	29 2���hz3���K� �rV�TRNDIAG.�LSw(:����� Ope��N� ~��nostic�����)VDEV�DAT�������Vis�D�evice�+IMG��./@/�/<�=k$Imagw/+7UP ES/�/?FRS:\?\=���Update?s List\?���� FLEXEV�EN��/�/�?����1 UIF Ev�O�O���,�t)�
PSRBWLD'.CMOϜG2#O�^?0�PS_ROB�OWELU���:G�IG�ϾO�?�O���GigE�(O��NߵA�)�AHADOW�O�O�Oi_���Shadow ?Change�����a�)RRCME�RRa_F_X_�_����PCFG Err{orq tail�_� MA�m�CMSGLIB�_�_�_`so�B6e��|0ico�+a�)_`ZD�O�o\o�o��ZDfPad�o l )RNOTI��o�ow���Notifiqc�� F�AG�� �՟����(���L� �p������5�ʏ܏ k� ���$�6�ŏZ�� ~������C�؟g��� ���2���V�h����� ���¯Q��u�
��� �@�ϯd�󯈿��)� ��M������ϧ�<� N�ݿr�ϖ�%ϣ��� [�����&ߵ�J��� n߀�ߤ�3�����i� �ߍ�"��/�X���|� ���A���e���� ��0���T�f����� ��=�����s���, >��b����'� K����:� Gp��#��Y �}/$/�H/�l/ ~//�/1/�/U/�/�/ �/ ?�/D?V?�/z?	? �?�???�?c?�?
O�? .O�?RO�?_O�OO�O ;O�O�OqO_�O*_<_ �O`_�O�_�_%_�_I_ �_m_�_o�_8o�_\o no�_�o!o�o�oWo�o {o"�oF�oj�o w�/�S��� ��B�T��x���� ��=�ҏa������,����$FILE_�FRSPRT  ��������A�MDO?NLY 1VU��� 
 �)�MD:_VDAEXTP.ZZZ3��䏻�ʛ6%�NO Back �file ���S�6)�����@�	� M�v�����)���Я_� �����*���N�ݯr� �����7�̿[�ٿ� ��&ϵ�J�\�뿀�� �϶�E���i���ߟ� 4���X���eߎ�߲� A�����w���0�B����f��ߊ��E�VI�SBCKs�]����*.VD����U��FR:\��ION?\DATA\��w��U�Vision VD��!�[� m����{��D����� z���3E��i�� �.�R��� �A�Rw� *��`��/� �O/�s/�/@/�/8/ �/\/�/?�/'?�/K? ]?�/�??�?4?F?�?�;�LUI_CON�FIG WU�����; $ �3x�{U�=OOOaOsO0�O�O�I%@|x�?�O �O�O__'\�OJ_\_ n_�_�_)_�_�_�_�_ �_o�_4oFoXojo|o �o%o�o�o�o�o�o �o0BTfx�! �������,� >�P�b�t�������� Ώ������(�:�L� ^�p��������ʟܟ ���$�6�H�Z�l� �������Ưدꯁ� � �2�D�V�h����� ����¿Կ�}�
�� .�@�R�d����ϚϬ� ������y���*�<� N�`��τߖߨߺ��� ��u���&�8�J��� [�������_��� ���"�4�F���j�|� ��������[����� 0B��fx�� ��W��, >�bt���� S��//(/:/� ^/p/�/�/�/=/�/�/ �/ ??$?�/H?Z?l? ~?�?�?9?�?�?�?�? O O�?DOVOhOzO�O �O5O�O�O�O�O
__ �O@_R_d_v_�_�_1_ �_�_�_�_oo�_<o@No`oro�o�o&h�`�x�o�c�$FLU�I_DATA �X����a�)a�dRES�ULT 2Y�e�p �T��/wizard/�guided/s�teps/Expert�o?Qcu ����������Skip G�pance an�d Finish? Setup�D� V�h�z�������ԏ����&h �`.�)`�e!�0 ��2`!��c�aA��ps������� ԟ���
��.�@�R� �2oy���������ӯ ���	��-�?�Q�)e@�)cA�3�E�W�g�rip*pu�ۿ��� �#�5�G�Y�k�}Ϗ� ��`����������� 1�C�U�g�yߋߝ�\� n����ߤ�b�g�%p�TimeUS/DST��?�Q�c�u����������
�?Enable��(� :�L�^�p���������P������ �b�a����������#�24 *������� 1C��y� ������	// -/?/Q/"4F\��$qRegion T/�/�/??+?=?O?�a?s?�?�?�AmericaϿ�?�? �?OO+O=OOOaOsO�O�O�)aym//�O��/�/#sditor �O7_I_[_m__�_�_�_�_�_�_� To�uch Pane�l  S (rec_ommenp)�_ >oPoboto�o�o�o�o�o�o�o�L��O�O5��O	_Racces �?����������,�>���Co�nnect to� Network M���������̏ޏ��@��&�8�J��H�^ !9+=S!_P�Introduct�/�����*�<� N�`�r������Ϻ�̯ ޯ���&�8�J�\�0n������� ��w������YVSafet�A$�6�H�Z�l�~� �Ϣϴ������ϩ��  �2�D�V�h�zߌߞ� ���������߷�ɿ� �[�k�}���� ����������1�C� �g�y����������������	-?[(�5��-�Q� ����"4F Xj|�M���� ��//0/B/T/f/ x/�/�/[m�/� ??,?>?P?b?t?�? �?�?�?�?�?��?O (O:OLO^OpO�O�O�O �O�O�O�O�/_�/3_ �/Z_l_~_�_�_�_�_ �_�_�_o o2oDoU_ hozo�o�o�o�o�o�o �o
.@�Oa#_ �G_������ �*�<�N�`�r����� Uo��̏ޏ����&� 8�J�\�n�����Q�� uן����"�4�F� X�j�|�������į֯ 诧���0�B�T�f� x���������ҿ俣� �ǟ)�;���b�tφ� �Ϫϼ��������� (�:���^�p߂ߔߦ� �������� ��$�6� ��?��c��Oϴ��� ������� �2�D�V� h�z���K߰������� ��
.@Rdv �G��k���� *<N`r�� ������//&/ 8/J/\/n/�/�/�/�/ �/�/����1?� X?j?|?�?�?�?�?�? �?�?OO0O�TOfO xO�O�O�O�O�O�O�O __,_>_�/?!?�_ E?�_�_�_�_�_oo (o:oLo^opo�oAO�o �o�o�o�o $6 HZl~�O_a_s_ ��_�� �2�D�V� h�z�������ԏ�o �
��.�@�R�d�v� ��������П⟡� �'��N�`�r����� ����̯ޯ���&� 8�I�\�n��������� ȿڿ����"�4�� U��y�;��ϲ����� ������0�B�T�f� xߊ�I����������� ��,�>�P�b�t�� Eϧ�i���Ϗ��� (�:�L�^�p������� �������� $6 HZl~���� ������/��V hz������ �
//./��R/d/v/ �/�/�/�/�/�/�/? ?*?�3W?�?C �?�?�?�?�?OO&O 8OJO\OnO�O?/�O�O �O�O�O�O_"_4_F_ X_j_|_;?�?_?�_�_ �?�_oo0oBoTofo xo�o�o�o�o�o�O�o ,>Pbt� �����_�_�_�_ %��_L�^�p������� ��ʏ܏� ��$��o H�Z�l�~�������Ɵ ؟���� �2��� �w�9�����¯ԯ� ��
��.�@�R�d�v� 5�������п���� �*�<�N�`�rτ�C� U�g��ϋ�����&� 8�J�\�n߀ߒߤ߶� �߇������"�4�F� X�j�|�������� ��������B�T�f� x��������������� ,=�Pbt� ������ (��I�m/��� ���� //$/6/ H/Z/l/~/=�/�/�/ �/�/�/? ?2?D?V? h?z?9�?]�?��? �?
OO.O@OROdOvO �O�O�O�O�O�/�O_ _*_<_N_`_r_�_�_ �_�_�_�?�_�?o#o �OJo\ono�o�o�o�o �o�o�o�o"�OF Xj|����� �����_'ooK� u�7o������ҏ��� ��,�>�P�b�t�3 ������Ο����� (�:�L�^�p�/�y�S� ��ǯ��� ��$�6� H�Z�l�~�������ƿ ������ �2�D�V� h�zόϞϰ��ρ��� �����ۯ@�R�d�v� �ߚ߬߾�������� �׿<�N�`�r��� �����������&� ����	�k�-ߒ����� ��������"4F Xj)����� ��0BTf x7�I�[����� //,/>/P/b/t/�/ �/�/�/{�/�/?? (?:?L?^?p?�?�?�? �?�?��?�O�6O HOZOlO~O�O�O�O�O �O�O�O_ _1OD_V_ h_z_�_�_�_�_�_�_ �_
oo�?=o�?ao#O �o�o�o�o�o�o�o *<N`r1_� �������&� 8�J�\�n�-o��Qo�� uow�����"�4�F� X�j�|�������ğ� �����0�B�T�f� x����������ᯣ� ��۟>�P�b�t��� ������ο���� ՟:�L�^�pςϔϦ� �������� ��ѯ� ��?�i�+��ߢߴ��� ������� �2�D�V� h�'ό��������� ��
��.�@�R�d�#� m�Gߑ���}����� *<N`r�� ��y���& 8J\n���� u�������/��4/F/ X/j/|/�/�/�/�/�/ �/�/?�0?B?T?f? x?�?�?�?�?�?�?�? OO���_O!/�O �O�O�O�O�O�O__ (_:_L_^_?�_�_�_ �_�_�_�_ oo$o6o HoZolo+O=OOO�osO �o�o�o 2DV hz���o_�� �
��.�@�R�d�v� ��������}oߏ�o� �o*�<�N�`�r����� ����̟ޟ���%� 8�J�\�n��������� ȯگ����Ϗ1�� U��|�������Ŀֿ �����0�B�T�f� %��ϜϮ��������� ��,�>�P�b�!��� E���i�k������� (�:�L�^�p���� ��w����� ��$�6� H�Z�l�~�������s� ��������2DV hz������ �
��.@Rdv �������/ ����3/]/�/�/ �/�/�/�/�/??&? 8?J?\?�?�?�?�? �?�?�?�?O"O4OFO XO/a/;/�O�Oq/�O �O�O__0_B_T_f_ x_�_�_�_m?�_�_�_ oo,o>oPoboto�o �o�oiO{O�O�O�O (:L^p��� ���� ��_$�6� H�Z�l�~�������Ə ؏�����o�o�oS� z�������ԟ� ��
��.�@�R��v� ��������Я���� �*�<�N�`��1�C� ��g�̿޿���&� 8�J�\�nπϒϤ�c� ���������"�4�F� X�j�|ߎߠ߲�q��� ���߹��0�B�T�f� x������������ ��,�>�P�b�t��� �������������� %��I�p��� ���� $6 HZ�~���� ���/ /2/D/V/ w/9�/]_/�/�/ �/
??.?@?R?d?v? �?�?�?k�?�?�?O O*O<ONO`OrO�O�O �Og/�O�/�O�O�?&_ 8_J_\_n_�_�_�_�_ �_�_�_�_�?"o4oFo Xojo|o�o�o�o�o�o �o�o�O_�O'Q_ x������� ��,�>�P�ot��� ������Ώ����� (�:�L�U/y��� eʟܟ� ��$�6� H�Z�l�~�����a�Ư د���� �2�D�V� h�z�����]�o����� �����.�@�R�d�v� �ϚϬϾ������ϳ� �*�<�N�`�r߄ߖ� �ߺ����������ӿ �G�	�n����� ���������"�4�F� �j�|����������� ����0BT� %�7�[����� ,>Pbt� �W�����// (/:/L/^/p/�/�/�/ e�/��/�?$?6? H?Z?l?~?�?�?�?�? �?�?�?? O2ODOVO hOzO�O�O�O�O�O�O �O�/_�/=_�/d_v_ �_�_�_�_�_�_�_o o*o<oNoOro�o�o �o�o�o�o�o& 8J	_k-_�Q_S �����"�4�F� X�j�|�����_oď֏ �����0�B�T�f� x�����[���� ���,�>�P�b�t��� ������ί�򯱏� (�:�L�^�p������� ��ʿܿ���џ� E��l�~ϐϢϴ��� ������� �2�D�� h�zߌߞ߰������� ��
��.�@���I�#� m��YϾ�������� �*�<�N�`�r����� Uߺ�������& 8J\n��Q�c� u�����"4F Xj|����� ���//0/B/T/f/ x/�/�/�/�/�/�/�/ ���;?�b?t?�? �?�?�?�?�?�?OO (O:O�^OpO�O�O�O �O�O�O�O __$_6_ H_??+?�_O?�_�_ �_�_�_o o2oDoVo hozo�oKO�o�o�o�o �o
.@Rdv ��Y_�}_��_� �*�<�N�`�r����� ����̏ޏ����&� 8�J�\�n��������� ȟڟ쟫��1�� X�j�|�������į֯ �����0�B��f� x���������ҿ��� ��,�>���_�!��� E�Gϼ��������� (�:�L�^�p߂ߔ�S� �������� ��$�6� H�Z�l�~��Oϱ�s� ������ �2�D�V� h�z������������� ��
.@Rdv ���������� ��9��`r�� �����//&/ 8/��\/n/�/�/�/�/ �/�/�/�/?"?4?� =a?�?M�?�?�? �?�?OO0OBOTOfO xO�OI/�O�O�O�O�O __,_>_P_b_t_�_ E?W?i?{?�_�?oo (o:oLo^opo�o�o�o �o�o�o�O $6 HZl~���� ���_�_�_/��_V� h�z�������ԏ� ��
��.��oR�d�v� ��������П���� �*�<������C� ����̯ޯ���&� 8�J�\�n���?����� ȿڿ����"�4�F� X�j�|ώ�M���q��� ������0�B�T�f� xߊߜ߮��������� ��,�>�P�b�t�� ������������ %���L�^�p������� �������� $6 ��Zl~���� ��� 2��S �w9�;���� �
//./@/R/d/v/ �/G�/�/�/�/�/? ?*?<?N?`?r?�?C �?g�?�?�/OO&O 8OJO\OnO�O�O�O�O �O�O�/�O_"_4_F_ X_j_|_�_�_�_�_�_ �?�?�?o-o�?Tofo xo�o�o�o�o�o�o�o ,�OPbt� �������� (��_1ooU��Ao�� ��ʏ܏� ��$�6� H�Z�l�~�=����Ɵ ؟���� �2�D�V� h�z�9�K�]�o�ѯ�� ��
��.�@�R�d�v� ��������п����� �*�<�N�`�rτϖ� �Ϻ����ϝ�����#� �J�\�n߀ߒߤ߶� ���������"��F� X�j�|�������� ������0����� u�7ߜ����������� ,>Pbt3� ������ (:L^p�A�� e����� //$/6/ H/Z/l/~/�/�/�/�/ �/��/? ?2?D?V? h?z?�?�?�?�?�?� �?�O�@OROdOvO �O�O�O�O�O�O�O_ _*_�/N_`_r_�_�_ �_�_�_�_�_oo&o �?Go	Oko-O/o�o�o �o�o�o�o"4F Xj|;_���� ����0�B�T�f� x�7o��[o��Ϗ��� ��,�>�P�b�t��� ������Ο���� (�:�L�^�p������� ��ʯ��ӏ����!�� H�Z�l�~�������ƿ ؿ���� �ߟD�V� h�zόϞϰ������� ��
��ۯ%���I�s� 5��߬߾�������� �*�<�N�`�r�1ϖ� �����������&� 8�J�\�n�-�?�Q�c� ��������"4F Xj|������ ��0BTf x��������� ��/��>/P/b/t/�/ �/�/�/�/�/�/?? �:?L?^?p?�?�?�? �?�?�?�? OO$O� �/iO+/�O�O�O�O �O�O�O_ _2_D_V_ h_'?y_�_�_�_�_�_ �_
oo.o@oRodovo 5O�oYO�o}O�o�o *<N`r�� ����o���&� 8�J�\�n��������� ȏ�o鏫o��o4�F� X�j�|�������ğ֟ ������B�T�f� x���������ү��� ��ُ;���_�!�#� ������ο���� (�:�L�^�p�/��Ϧ� �������� ��$�6� H�Z�l�+���O����� ������� �2�D�V� h�z��������� ��
��.�@�R�d�v� ��������}��ߡ��� ��<N`r�� ������� 8J\n���� ����/���� =/g/)�/�/�/�/�/ �/�/??0?B?T?f? %�?�?�?�?�?�?�? OO,O>OPObO!/3/ E/W/�O{/�O�O__ (_:_L_^_p_�_�_�_ �_w?�_�_ oo$o6o HoZolo~o�o�o�o�o �O�O�O�O2DV hz������ �
��_.�@�R�d�v� ��������Џ��� ��o�o�o]����� ����̟ޟ���&� 8�J�\��m������� ȯگ����"�4�F� X�j�)���M���q�ֿ �����0�B�T�f� xϊϜϮ���ѿ���� ��,�>�P�b�t߆� �ߪ߼�{��ߟ��ÿ (�:�L�^�p���� �������� ����6� H�Z�l�~��������� ��������/��S ������� �
.@Rd#� �������/ /*/</N/`/�/C �/�/{�/�/??&? 8?J?\?n?�?�?�?�? u�?�?�?O"O4OFO XOjO|O�O�O�Oq/�/ �/�O	_�/0_B_T_f_ x_�_�_�_�_�_�_�_ o�?,o>oPoboto�o �o�o�o�o�o�o�O _�O1[_��� ���� ��$�6� H�Z�o~�������Ə ؏���� �2�D�V� '9K��oԟ� ��
��.�@�R�d�v� ������k�Я���� �*�<�N�`�r����� ����y���������&� 8�J�\�nπϒϤ϶� �������Ͻ�"�4�F� X�j�|ߎߠ߲����� �����˿ݿ�Q�� x������������ ��,�>�P��a��� ������������ (:L^�A� e���� $6 HZl~���� ���/ /2/D/V/ h/z/�/�/�/o�/� �/�?.?@?R?d?v? �?�?�?�?�?�?�?O �*O<ONO`OrO�O�O �O�O�O�O�O_�/#_ �/G_	?_�_�_�_�_ �_�_�_�_o"o4oFo XoO|o�o�o�o�o�o �o�o0BT_ u7_��oo��� ��,�>�P�b�t��� ����ioΏ����� (�:�L�^�p������� e��ӟ���$�6� H�Z�l�~�������Ư د����� �2�D�V� h�z�������¿Կ� �����۟%�O��v� �ϚϬϾ�������� �*�<�N��r߄ߖ� �ߺ���������&� 8�J�	��-�?ϡ�c� ���������"�4�F� X�j�|�����_����� ����0BTf x���m�������$FMR2_�GRP 1Z��� ��C4  B��	� ��;M8E�� F@ cǂ5Wo�
8J���NJk�I'�PKHu��IP��sF!��{?ǀ  ��89��<9�8�96C'6<�,5��{Ag�  /+BH5�B�10 !@�3]3;"�33�7x]/n-8@UUT�*�@9 � {��>u.��>*��<����{>���>���l=<��=��U�=�v!>1�
{:�ܜ:�2B8'Ŭ9�IR7���9f�͛/$?o/!?Z?�E?~?i?�?��_C�FG [T ��?�? OO�;N�O 
F�0HA M@�<RM_�CHKTYP  ���&(� R{OMc@_MINi@������@�T X�SSB�3\�? 9�O���C�O�O�5TP__DEF_Oz���&	WIRCOM�h@_�$GENO�VRD_DO�F���G]THR�F dzdUdMT_ENB9_{ MPRAVCu]�G�@ �[�F@ G��@�GAw\H͊#Iv0�Iά �?�Oo�o(oK*� �QOUc�PAKRK<�@��oIo�o�o��o��C�  D��o�h1A|A$ B��L.rN�i�O�PSMTd�Y*�@t�$HOSTC�2s1e�@����7 MC��T{����  27�.02�1�  e�_�q�������M��Ə؏��������	�anonymous#�Q�c�u��������6������� F�'�9�K�]�o����� ����ɯ쟆�0��#� 5�G�Y�k�����ҟ�� �׿�����1��� �g�yϋϝ������ ����	��-�p��ϔ� ���ߺ�ܿ�������� �H�)�;�M�_�q�� ���Ϲ��������D� V�h�z�|�R��ߑ��� ���������!3 Eh������� ��*�<�N�PA�� ew������� �//<n3/a/s/ �/�/�/���/$/ ?X9?K?]?o?�?� �?�?�?�?�/�?B/#O 5OGOYOkO}O�/�/�/ �O�?�O,?__1_C_ �?g_y_�_�_�_�OT_ O�_	oo-o?o�~�q�ENT 1f�y��  P!�_�o  �p~o�o�o�o �o�o'�o3\ �D�h���� ���G�
�k�.��� R���v���鏬��Џ 1��U��N���z��� r�ӟ�������ޟ,� Q��u�8���\����� ᯤ����گ;���_��"�QUICC0 l�H�Z���~�1�������~�2����[��!ROUTER�\�8�Jϫ�!PC�JOG�χ�!�192.168.�0.10��z�CA�MPRT����!b��1��#�
�RTu��'�9ߚ� !So�ftware O�perator Panelw������`dNAME !~mj!ROBO����S_CFG 1�emi ��Auto-st�arted�DFTP�O���O�_�� �O��������c_>� P�b�t����+����� �����@\�n�� a����x���� ��'9Kn� �������O�O �O�OV,/�k/}/�/ �/�/v�/�/�/?? B/�/U?g?y?�?�?�? �//(/*?O^/?O QOcOuO�OJ?�O�O�O �O�OO�O)_;_M___ q_�_�?�?�?�_�O�_ 2Oo%o7oIo[o_o �o�o�o�_�olo�o !3EW�_�_�_� �o�o�����o A�S�e�w����.��� я�����\n� �s��������͟ߟ 񟴏�'�9�K�]��� �������ɯۯ�0� B�T�f�h�Y���}��� ����ſ������� 1�T�ֿg�yϋϝϯ������_ERR �g�����PDUS_IZ  V�^t�����>	�WRD� ?J�7�� � guestV�I�[�m�ߑߣ����SCDMNGR�P 2hJ����7�V�8V��K�� 	P01�.03 8� �  e�?���  ;  ��  � ��������@��-�������x����0���y� d����,�>�P������  	D��d����������_GROU��i*������	���]5{�QUP�3��������TYC �����TTP_A�UTH 1j��� <!iPen'dan��%`Ϗ��!KAREL�:*%.@KC�UewM VISION SET����V�K�� J(@:�^p�����CTRL� k����%V�
�D�KFFF9�E3�5�FRS�:DEFAULT�3,FANUC� Web Server3*! 5���1� C���/�/�/�/�/?���WR_CONF�IG l�� �3/��IDL_C_PU_PCR V�sB�8�u0 BH[5�MINf<!�y5GNR_IO���V����]0NPT_SIM�_DO�6�;STAL_SCRN�6� ���INTPM?ODNTOL�7�;�!RTY�8u1�6� N��ENB�7��Y4OLNK 1m��E�}O�O�O�O�O�O|�OaBMASTE�0���aBSLAVE �n��URAMCOACHE_�2O��O_CFGI_`CaS�UO��l_]RCMT�_OPR �2�ʟSY�CLH_{UL _AS�G 1o��#�
 �Oo o2oDoVoho zo�o�o�o�o�o�o�o\�K�RNUM����
]RIPF_XWRTRY_CN�_{U�1(���|A��� ]R�PfRp'^=з=�]0�P_MEMBER�S 2q��� $�%�r����w���]0RCA_AC�C 2r��  �V�# 
�3� /� 3y O 5��(�� S��5`�H�c�U� � V�5�BUF�001 2s��=� �u0  ou0�փބ�ބ#ބ(V�� 	�փ

���+�;�L�[��m�|�������������Z��փ~�~�U!~�1~�B~�Q~��c~�r~��u0(� M�u0��`x�u0I_�+��~��~���u0�s8}րuփ�,��Cu0$�QYu04��@�%?�  o?�4փE&��T&�=�6�>p�E� r0��ք ք/ք��V��bքqք�քU�ք�ք�ք�ք	�փ��2��҃ց܁�ց������k(
��ց���� ��%��-��5�� =��E��M��U�� ]��e��m��u�� }�ց������������ ���������������� ����Ő��͐��Ր�� ݐ��吉��ց���� �����������ցx��$�_@�,��!�5�!�F�D�t(L�N�T��]��e� ᢮�t��}�ᢅ����q�`��ᢝ� ᢥ�᢭�ᢵ�ց��3ɯ҅�^"��^" ��` ��8���"� #�"%�3�"5�C�" E�S�"U�c�"e�s� "u���&񄓓��ҕ� ���ҥ����ҵ�ó�� Ő��͐��Ր��ݒ� ���&�������� ���&��+�*�-� ;�*�O�D��M�[��� ]�k��·�t����� �������¥�����X����gQ2t��4,%&�&�<&�K���25�HIS��v�� �S� 2�023-07-2���Y"{O�q8 U�p����������������V�Y&E�19Q�|B;��p:m�L^p���p����s!8Q�,>Pbtd�Y!�Y!׀���ҫ�s!�:�s
��7��q� /"/4/F/X/j/|/�/ �/���/�/�/?? 0?B?T?f?x?�/�/�? �?�?�?�?OO,O>O PO�?�?�O�O�O�O�O �O�O__(_z#�ȠP/�A�e�:- dU��Qc3_�_�_�_�_�_�oo1>  dA �d0oo�o�o�o �o�o�o�o��|_E�Wi{���� �c�io��r�- ' L�z�^iO{O �/�A�S�e�w����� ����eO�����+� =�O�a�s�����Ώ�� ��ߟ���'�9�K� ]�o�����ʟ��ɯۯ ����#�5�G�5_"� ��T_f_0e�ӹ� ƿؿ���� �2�D�h2oDoVh"� U� �ϲ����������� 0���f�xߊߜ߮� ���ߛ- ��߼-  �- �����B�T� f�x���������� �-��,�>�P�b�t� ������������� (:L^p�� �������� $�6HZlZ�l�I_�CFG 2wz�� H
Cycl�e Time��Busy�Idyl��min}=�Up���Read�gDow�� �}�Count��	Num ���ȩ`,S�7!EQPR�OG�xz����p/�/�/�/�/�/�?�@USDT_ISOLC  z����pJ23_�DSP_ENB � B;�c0INC� ys=S�P0A �  ?�  =�?��<#�
O1�9:�o �1�?�?�S��?O\7OB� C�l3��6"AG_GROUP 1zB;;�r<� �3(�	nOO?��/�OS�Q�O�O�O_�O0_�B_T_f_��?IG�_IN_AUTO�/D�:c0POSRE�*O<FKANJI_�MASK�V�ZKA�RELMON {z�h/S�y+_DoVo@hozo�o�b�#|�'�~3S��e�_4K�CL_L�PNUM�p0�o$KEYLO�GGING�`����q{5� LANGU�AGE z��Jp�DEFA�ULT Xqh�LGf�}�*��Sѽx�0�  R��H  �S�'�� + �SЛS�?)7�;��
�q(U�T1:\�o�  ����0�=�O�a�x�������(3o�c��LN_DISP �~�?��O�O��O�CTOL9�S�Dz�� K1�1O�GBOO	Kq0i}d���������X�|����ϟៀ���us�'��	m��yjA%;o�?�1�k�_BUFF 2��B; �S�2 �����*2ү�� � -�$�6�c�Z�l����� ��Ͽƿؿ���)� ��2�_π3��DCS ��)�2�1$�c������������v�IOw 2��� �3�jA�6�F�X�j� ~ߎߠ߲��������� ��0�B�V�f�x�������������ER/_ITM?>d�_?� Q�c�u����������� ����);M_�q���I��SE�V�`s=�TYP?>.�!3��Q�RSTt�SCRN_FL 2��� ��ϧ���0�//DTPp??��C�NGNAMpl4��Jrr�UPS�SGI\�U{5�!�_LOAD'@G �%@*%DMA�Yɥ�/G�MAXU�ALRM�b�QC���{5
�"�!_PRD�$�P a�%�� C��i�ٯè)3H@�P 2�w� �ZƦ	O!t�0��0�P?���2�?�?�?�? ���?+OOOO2ODO�O pO�O�O�O�O�O_�O '_
__]_H_�_l_�_ �_�_�_�_�_�_�_5o  oYoDo}o�oro�o�o �o�o�o�o1U gJ�v���� �	��-�?�"�c�N� ��j�|������̏� ���;�&�_�B�T��� ������ݟ�ҟ����7��'DBGDEF �25?1>1@�R��_LDXDISA�m ?+�MEMO_{APg E ?@+
 d����ү������,�>�� F�RQ_CFG ��27h�A �@i���!�<?4d%A�Э�R�d�z2�2;��4*��/�� **:�!��� ȟ�!�,�>�k�b�t� �ϘϪ���#�25 ���`��'�� �6�,(�� ~���lߩߐ��ߴ��� ���'��K�]�D���h�������*IS�C 1�@)� � )�#��4i�9�$�r�]��������_MSTR� ����SCD 1�������� ,P;t_q� �����& L7p[��� ���/�6/!/Z/ E/~/i/�/�/�/�/�/ �/�/ ??D?/?A?z? e?�?�?�?�?�?�?�? OO@O+OdOOO�OsO �O�O�O�O�O_�O*_ _N_9_^_�_o_�_�_��_�_�_�_o��MK�g������&o$M�LTARMf��:۷Qb �b���o�dQ�METPU܋�b����ND�SP_ADCOLx�ef��nCMNT�o �eFN�`�o�gFSTLIw�� ���g~�c��|�t�ePOSCF5w=�nPRPM�o�y�ST�`1��� 4��#�
��� �!��!�#�5�w�Y� k��������ŏ׏� ���O�1�C���o��a�SING_CHK�  $MODAe���OkQn���DEV 	��	�MC:�HSI�ZE��`ȿ�TA�SK %��%$�12345678�9 `�r���TRI�G 1��� l Q�����Lٮ��L�B��YP-�L�Ք��E�M_INF 1��ۻ`)AT?&FV0E0��k��)S�E0V1&�A3&B1&D2�&S0&C1S0}=Z�)ATZk�����Hÿ�z�߯���A�C���g�Nϋ��� Q���u������� �Ͽ@�w�d�v�)Ϛ� U߾��߷��ߧϹ�*� �����r�}�7ߨ��� �������&��J� \���3�E�W�i��� ����5�4��X |�u�e�w���� ����0B��f�� EO�{��// �>/�'�/K �/�//�/�?�/'?�L?3?p?�NITO�RPpG ?�  � 	EXEC�1c�22�83�84��85�8���67�88
�89c�2:"D�2 D�2D�2D�2D�2 D�2D BDBDB�C2%H21H2=H2�IH2UH2aH2mH2�yH2�H2�H3%H3�1H3�2��R_GRP_SV 1�@�� (w���<�� ��>%���6����u�=���J�_D�20�ySION_D�Bɐ�͝a  ��`�☾T �Z`��W��pr�>f0N   #v�W�G�-ud1��/oAoSo�aPL_NAME !Q��|`�!Def�ault Per�sonality� (from FsD)�P�bRR27Q� 1�L�XL��x|a�P dzr�o�o�o�o# 5GYk}��� ������1�C���2�on���������@ȏڏ������<]� :�L�^�p���������@ʟܟ� �[i*�)�":�
)�^�]dPM��� ������ү����� ,�>�P�b�t�����g� y�ο����(�:� L�^�pςϔϦϸ��� �ϫ����$�6�H�Z� l�~ߐߢߴ����������� �2� F�@ G&h G�]gSP  �_�q�]bd[�C���� ������D�7�Zj��	�p��=�@� -� X�N�`�r����������SP�0��	]b-�	�`B�<N`:�oA�b����? A�  �	W�kV]`�S ]`�PCT��s � h�`)  �  u$�T &"�C�gyd���\kR6R 1��ti�P*0 �� f2|`  @oD�  !?�#X,?]`!]a�A/��%iJ-;��	l,"	 ��pJn �NP`e  � �� � �� � ���"SPK�K� ��K=*�J����J���J9٧�U�p��/�SP@_f��"j�@�(E14!�/��#�N����;�f,1�� �a�������-�@·�  T1�HZ0�Z0� �/  >c��=��>�]a�ǿ����l? �?�2-!�3�&.W p�Pm P� }��P�  ��P��F�*O�%	'�� � HBI� �  ����&:�ÈlOÈ�=��̈́E�"@�O�@�>!�O/K"���&&�&�Q_ � '`.T�!-0@2?��@����"=0�@A?C� C�PC��� Ca0Ce0C�i=%��A�%� 0 �Pl~�-hhX�'B�P�Q���A�U]aDz�on?3ooCo io�O�dIA�R�TZ��A����  �4@?�ff���o�onoC  #{�!8�@9Gz>L�@�0(!�*(�@uu�0�v�i{!t#�t$�C?]t�@,��<�
6b<߈;�܍�<�ê<���<�^¬/d�C�A�K"�#|,"� ?fff?�@�?&&���@�.�8��J<?�\�D�N\��I�R!�-$ �)%|�'��
�`$�o Џ���ߏ��<�'��`�r�]����He�F | ��ҟ����m������J��F�  F����BG�d GC�qV���R���ů�� �ԯ���1��U�@� �O���F�IG/�ӿ1����m��0�B�T�:��o�{�33ϩ��@�ϸ������{An� ��_�EC��U��ϲ�d�?�؃ߊ��ߴ���I�i4����C CfPa0�¸���0؜�@�@I����B>�)A�C��AIA���@�?\����ú�@ �������=q�A��Ay�I3�3@0��@���C�1�������(��C���b��=q�Ů�����H�� G�� �G�B�I��(?E�� C�e�� �I"L�J��HV@G5� �E�x C��I�3�J0�G���I�� 0 C='�߀�k����� ����������"F 1jUg���� ���0B-f Q�u����� /�,//P/;/t/_/ �/�/�/�/�/�/�/? ?:?%?7?p?[?�?? �?�?�?�? OO�?6O !OZOEO~OiO�O�O�O �O�O�O�O __D_/_ h_z_e_�_�_�_�_�_:y�(������r���$e�U��xo&o9�3�8�@o<Ro9�4Mgulo~o�9ѴVwQ�o�o4p�+4�]�m �i�o(L:|u�%P�rP~~�������_�����{R���G�2�W�}�h�  �`��ˏ��� ڏ����F�4�j�X�p�z��������ԟz����4�"�X��F�|���  2 wF@9�G&h����9�B�&��)�&�C�&�9�@-��9�o�+�=�O��� ����Ħ�GAw�\]�����ɿ7�?���|p9�t�9��9���{�
  ֿ9�K�]�oρϓϥ� �����������#�z�����hk�y���$MR_CAB�LE 2�hx� �ћqT�p	@����?>𦡆т�K��кƠ��C���ޱO8�tB��]��8��ް.ޱ�F\!�޶�ߕ���>��š��C�N��|�����a}9`r���	P��e�����L  ���C�֠:������^�a��!ްޱOE� "�4��ՠ��y�By�ԡ��HEو��ls�޵;�aZv�/ߘ���k�� ����C��L�>�8�f� \�n�������������P?��H�� oq< ���ܸ����ܸ*,** �\�OM �i������ Ël%�% 234567O8901i{ fH��ް�ް�ް�ޱ
�n�ot sent �5�WpuT�ESTFECSA�LG#�egۺ�d�.$��
>$����p޴�޷Y/k/}/��/ 9UD1:�\mainten�ances.xm�l�/�/  ���DEFAUL�Ta�\�GRP 2=�M  pė��޵  �%1s�t mechan�ical che�ck�ޱ�z3鰄1�?��[ph��?��?�?�?�?޲R3co�ntroller b4,O{?PO���?|O`�O�O�O�OAMY=,�O޲"8SްQ_��kG8_J_\_n_�_�JCO�__�_�6/_oo(o:oLoB�C[0geW2. b?atteryPo�_�o��	�_�o�o�o�o�_i@dui@awble  D50 Pq��`���o������Addg�reas;޷f�B�-ް�#���{@P�b�t�����A
dd�oi�/��+��?��&�8�J�\�AXdj7޶����<ް������
�؟���� �#|too�����>ǟ������ү�A�Overhaul�Ow��"� xް,�3�:5��`�r�������ް$Q�пSV�� O�$�6�H�Z�l� ����߿�Ϲ����� � �2߁�VߥϷ��� �߰�������5ߝ�� k���d�v���� ������1��U�*�<� N�`�r���������� ���&8��\ ����������� �M"q�X�| �����7I /mB/T/f/x/�/� �/�/�/3/??,? >?P?�/t?�/�/�/�? �?�?�?OOe?:O�? �?�?�O�O�O�O�OO �O _OO�OsOH_Z_l_ ~_�_�O�_�__�_9_ o o2oDoVo�_zo�_ �_�o�_�o�o�o
 ko@�o�ov�o�� ���1�Ug<� �`�r��������̏ �-��Q�&�8�J�\� n�������ȟ�� ���"�4���X����� ˟����į֯���I� �m����f�x�����p����5��	 T¿ ���*�4�F�X�j� |ώϠϲ��������� ��0�B�T�f�xߊ� �߮����������� ,�>�P�b�t����޼�  �b�?�w  @�  � ��	�����H�Z�l���*��**  @�>�7����������p,>��e� ^���A���u� ��EWi�Ug y�����/ �/-/?/�/u/�/ �/��/�/�/??��/;?M?_?�/�/����$MR_HI_ST 2�>��0�� 
 \
�$ �23456789C01�?�4�?���?9�)O;O�?$O��O �O�O^OpO�O�O_�O �O_I_[___6_�_ �_l_�_�_�_o�_3o �_Woio o�oDo�o�o zo�o�o�oA�d��0SKCFMAPw  >��0)8�1�`IYu�ONREL  ƚ5rq�0[rEX_CFENB�w
ps�Xu�qFNC��tJOGOVLIM�wqd�3�[rKEY�w���_PANp�x+�'�[rRUN ��,�SFSPDT�YP�x�uZsSIG�N��tT1MOT���q[r_CE_�GRP 1�>�rs�2ڰ9���c�� 8��8&�g����B��� ��x�埜�ڟ�ҟ?� Q��u�,�����b�ϯ ��ȯ���)�;�"�_�������|����7[qQ?Z_EDIT��lw���TCOM_CF/G 1�h}�u��&�8� 
��_AR�C_�r�5�yT_MN_MODE�����yUAP_C�PL]��tNOCH�ECK ?h{ @ ������ ��,�>�P�b�t߆���ߪ߼����ߍ{NO_WAIT_L��l�ՀNT���h{�w��c2�_ERR&߁2�hy�1�6��� ���*��q�����w��O`�g�| 
��;��0��a<O�00 ?�5�O�5��p"�Y�_PARAMa�h{��� ������1�� = O0 8ZlHx��`��������.��R��ODRD�SP\ã��xOFFSET_CARజbψDIS��S;_Aw�ARK����OPEN_FIL�E���;��S�OPTION_IO!��3� M_PRG ;%hz%$*E/W.��WO������00�%�d.2 ; p	  �d� �C�#��h�!�f����hRG_D?SBL  �7rq�K�?eRIEN�TTO�p�aC��pqqA� hUT__SIM_D'or���hVlLCT �<�粛$;��9�e=d`7_PEX��n�4RAT� d�u��4�UP �q>�{ �OOO�BOPI�$��2ރ��L�XL�x[3�0C�O�O �O�O�O�O__(_:_ L_^_p_�_�_�_�_�_�_�_ o�g2�O/oAo Soeowo�o�o�o�o�o B�o�o1CU gy�������f��o�~9@�!�N�P �K�]�o��������� ɏۏ����#�5�G� Y�(�:�������şן �����1�C�U�g� y�����l�~�ӯ��� 	��-�?�Q�c�u��� ������Ͽ�s�¯��C� �2͠4AP� b�Gυϓ���A�����ϭ������� !�3�Q�W�uߗ���{ 0��������	`���x�!�x�:�o@1�?�Q�c�u�A�S  ��V+��!�+�21� 9����s  h�p �)  �  u$�����)��&�@_�J���^fBl@O�0�1����� {D��0 ��$  �� @D��  ��?����X,?+���+�D��������  �;�	l��	 ���pJ�3 �����*  Կ � � �I �� �Ou�H(���H3k7HSM5�G�22G���GN�3h��(ϙL�u�CH50�R50������r�û��׾  ��� ��� �)��m�AK��µ+�²g���801 i�o��u����� Up m3�P00� _�  � ���u��q�	'� �� "I� ��  ���o�=����1/C+�@Y/_ Z�!�/��"!�����q�NA0�/�  'R0�$���CNA0C���*C.p ??�q�p�Az
�b0lwhhXn�B� �1��~�p!�5��zn��?3 �?�?O.OU/GD!N2�K4a+���>�@?�ff�ϏO�O3O ���O�KA18+��OZ>LS ���J(+�:U�EV^I�@99�#?"T� ,�A<
6b<���;܍�<����<���<�^��q�_�AAp+����#���?fff�?p ?&�PD@��.�R�J<?�;\�	bN\��U2 �Q�@��Ao��`o�W %�O�o�o�o�o�o�o �o%7"[mD �|�,oNoPo����xF�  F��~+�G�d GCFQ �T��d���u����� ҏ��������/M� �&
������2� ������J��O�[�3pޟw�b�������
<�A3�墚?+��C�����w�)�?Ƀ�H�O���s�
Ķ4�ț�C��C�࿇�b��b�a���@I�	B>��)A�C�AI���A��@�υ?\������ú@ �������=q+��R!>�I33@0���@��C�1����[�������C��'���=q�Ů���	H�� �G�� G�B��I��(E�� �C�^l��I"L��J�HV@�G5� E�x �C���I3�J�0�G���I��� E@� C ��E�0�i�Tߍߟ� ���߮��������/� �,�e�P��t��� ��������+��O� :�s�^����������� ���� 9$]o Z�~����� ��5 YD}h �������/ 
/C/./g/R/d/�/�/ �/�/�/�/	?�/-???�*?c?N?�?r?�?>�(�I���^opR��<�5�5���?�?@�3�8�OO@��4Mgu1OCO@���VwQ]OoO4p�+4�]�M�I�O@�O�O�O_�L:�P�R	PC^>�_�l_�?x_0�_�_�_�[R�_�_`o�_oBo-o  �@�EoWo�o{o�o�o�o�_Q��o/{ 5?uc���?�������A��O�  2 F�@@�G&hl����@�B����ձC	��@�@򯷏ɏۏ ����"�@��oL�`^�p�����@�?���TAP@��d@�@�r<���@�
 �� ���"�4�F�X�j�|� ������į֯�?ʶ����-K�y���$PARAM_M�ENU ?�E��  �DEFPUL�SE��	WAI�TTMOUTL��RCV_� S�HELL_WRK�.$CUR_ST�YLJ���OP9T����PTB�����C��R_DECSNW�4U���%�N� I�[�mϖϑϣϵ����������&�!�SSR�EL_ID  �E]Q�5�USE_PROG %0�q%"߇�6�CCRc��G�]Q8���_HOSoT !0�!���ߔ�TTP���ӿ������4��_TIM�Ea�G֯�!�GD�EBUGE�0�6�G�INP_FLMS�K]��T�P���P+GA�� |�;����CH���TYPE
-�9�!��Q�z� u�������������
 )RM_q� ������* %7Irm�����/��WOR�D ?	0�
 �	PRy��SMsAI���RSUͱ�=#TE��S�	��J"COL�Uf)�/Z��Lc� �@��`�ȯ�dq�TRACECTL 1��E�:� AP%/ &'AP;P�.��&DT Q��E�0� D � �;�+0̐10�[Q92��92Ԑ92.3��56Ȑ12f5/4�/4	/4
/4/4�/2�=4�E4�M4��-4�54�e6/4�/4/4G�12/4�/4/2� D�DTp	B��	B!D"�D#D$/13S���4��4�=4��E4�M4�-4�54��e4��4��4��4�N�4� DED�DD�12>3�E4�M4,?>?P?b?t? �?�?�?�?�?�?�?O��OC��	BWDS�BT�T�!XC�S�TU�T�T��D�-f(�E�EFS�MT�UT0! XCVOhOzO�O�O�O�_ �O�O�O
__._@_R_ d_v_�_�_�_�_�_�o �_oo*o<oNo`oro �o�o�o�o�o�o� &z'1KEo������� ��ɟ۟����#�5� G�Y�k�}�������ů ׯ�����1�C�U� g�y���������ӿ� ��	��-�?�Q�c�u� �ϙϫϽ�������� �)�;�M�_�q߃ߕ� �߹���������%� 7�I�[�m����� ���������!�3�E� W�i�{�����k����� ����%7I[ m������ �!3EWi{ �������/ ///A/S/e/w/�/�/ �/�/�/�/�/??+? =?O?a?s?�?�?�?�? �?�?�?OO'O9OKO ]OoO�O�O�O�O�O�O �O�O_#_5_G_Y_k_ }_�_�_�_�_�_���_ oo1oCoUogoyo�o �o�o�o�o�o�o	 -?Qcu��� ������)�;� M�_�q���������ˏ ݏ���%�7�I�[� m��������ǟٟ� ���!�3�E�W�i�{� ������ïկ���� �/�A�S�e�w����� ����ѿ�����#���$PGTRACELEN  "��  ���!��7�_UP �����f��n�R�g�7�_C�FG �f�TP�!�g������ϸ�I���  ����{�DEFSP/D ��� �I���7�H_CON?FIG �f�N�W !�!�d-�M�F�  �0�P�����L�!��7�IN~~�TRL ��Ͳ��8��a�PE����f���,�\��7�LIDù���	��LLB 1��� �M�B�<�B4�� �M�%��Pպ� <o< �?�O� n�O�f������� ���"���<�j�P�r�����8������� 
Q�@3Ev�ٿGRP 1�����"�@��
����!�AM�D��@ D�@ C5f� @ �1���0�	�	,�,����uG���´F(BIpP:L�p��!�>�l7>�ú��/.� =�-=%�T/ Q//N/�/r/�/�/0/��/�/�/?)??  #DzN3W?!�
>?? .?�?�?�?�?�?�?�? !OOEO0OBO{OfO�O�O�O�J)�A
V�7.10beta�1�� A��=� R�!�A!��@�?!G�Q=y��#�B���$Q@�����B�l�4Q@�A���QT� �Oi_{_�_�_FTp���<��_�_�_�_ .� ��O��O�0oBo@,ofoPo�o�A-�p��u0�mf��o��o���@�AWP�R�c� B��B�>0uB�Hfs�d!�!�LPuM���d����r
�cx�tx��h��$|�����0��<�-�@�F�0�A��33`�������KNOW_M  ��"�����SV ��C�]�m? �� $��oH�3�E�~�!�����M��� �jR	��ѐlb���^���hhXd��1q� (�0u�8�4�����MR�� ���&�oj3�������OADBANFW�D����ST�1 k1�f��4�� �Y�!

��.�_�R� d�v��������п� '���]�<�Nϓ�r�@���ϨϺ����2��8��	�ݠ�<3�߂�3�/�A�S��4 p߂ߔߦ��5���������6�(�:�L��7i�{����8`���������MA֠���b�OVL/D  ��~��PARNUM � �������SC-Ha� o�
����8	�UPD�����#bb�_CMP_0��d����'�z�ER_CHK�����˒���RqSu�ٯ��_MO֯��_�a�_RES+_G����
V_�� ch������ �/
/;/./_/R/d/7�DT�/9o� �/�/�/;���/?? ;�!?@?E?;h�`? ?�?;���?�?�?;���?�?O;V 1���vߠ��@`}�\�THR_IN�Ru�f��dqFM�ASS~O Z�GM�N}O�CMON_QUEUE �����
�Qa�N U��N�F�H SEND8Q#YEXE._U�D BE-P_ SOP�TIOW,PPR�OGRAM %��J%P<O��RT�ASK_Ic�u^O?CFG ��O����_
`DATA���&kP�
2ʕyo �o�o�o�olo�o�o	 -�oQcu�:o�INFO���Wm� �DC����(�:� L�^�p���������ʏ ܏� ��$�6�H��w�t�Wl r)	a��K_a�i�~���ENBd�ѹ�2�ԘGa2̙�� X,		�=���� ���@�N�9�$��8�8�`D���_EDIT ��o����dWER�FLOXdC�RGA�DJ �}�A����?
���AϦQ�������??�  Bz��ga<8�
�v%$�\�è�r-�g�2���r	�H�@locBB=P���q@'�ǽ�*۰/ݲ *�*:�ֿ��q<��.@A��ſ�@K�@�c���\I)#����1�[ϩ�g�������w�A.@u����� ��O���K�5�/�A߻� e߷ߡߛ߭�'���#� ����=��y�s� �������������k� �g�Q�K�]������� ������C��?)# 5�Y���� ���1� mgy����� �_/	/[/E/?/Q/�/ u/�/�/�/�/7?�/3? ??)?�?M?�?�?�?�?{�	&o0OŠOWOBD�t$ qO�KEO�OAO�O�O	�PREOF ��ŠŠ�
ϥIORITY�W���ӡMPDSaP�Q��A�7WUT�V|��ΦODUCT�Q�}��O��OGg�_TG���R��vR�HIBIT_DO����[TOENT �1�}� (!?AF_INEaPo~g!tcpo>Gm!ud6oon?!icm^o��vRXY��}��š)� ��o�oŠ��o�e�o:! ^EW�{���@����6�H�*uS���A�J�����£�>Ԥ�Ѷ�/���z��¤�r�}�A~;�,  �P�}�8�J�\�n�ť�߆Zߏ����ҟ�£�]�ENHANCOE �i�}�A�AdޏD�+�rV�D� _�SɡӡPORT�_NUMbSŠ�.Uӡ_CART�RE���l	�SK�STAaW�[SLGmS`ٸk�;��HPUnothingL�)�;�M�]����������_�TEM�P څY���5�q�_a_seiban�OϯO(�N�9� r�]ϖρϺϥ����� �����8�#�\�G߀� kߐ߶ߡ��������� "��F�1�C�|�g�� ������������	� B�-�f�Q���u����� ��������,P ;`�q����������VER�SI@P�WQ �disable�^���SAVE �ۅZ	2670/H769'��!4���po� 	�	(kR�?;+2/ESe@O/x/�/�/�/�*g,���/z�n_�P 1ܸk�20
B�5�<?N?�7�@URGEb�B�P�^�aWFz0�QdT�pVW`�4LQ���WRUP_DE?LAY ݼ��5�R_HOT %�FnQ3�O�5R_NORMAL�8�R
O<_O.GSEMI>OdO|�O�AQSKIP3	�p�+3x�O_ _0_�M�5W_eWO_�_ �_�_o_�_�_�_oo 'o�_Ko9ooo�o�oYo �o�o�o�o�o�o5 #Ek}�U�� �����1��U��g�y��5�$RBT�IF�4��RCVT�MOUէå����DCR3��I� ��AC�}��C���C����?���>�9��<<�Mä��`��2	1��$,��� ��(9��OC�?_ �<
6b<߈�;܍�>u.��>*��<����U���?�����  ��ߟ���'�9�K��]�o��������ERD�IO_TYPE � !=����EDP�ROT_CFG ���G�4BHf3E���A2��7 ���B� �T� b�����:�����п�� c�ϐO(�G_I�;�Y� [�mϣϑ��ϵ����� �ߡ���E�3�i�W� ��{ߝߟ߱���	�� -�/���?�e�S��w� ������������+� ��O�=�s�a������� �����������K 9o]������ ���5#EG Y�}����� /�1//U/C/y/g/��/���/����INOT 2��9J��ǱG;� ?&;s���<N?�f�0 l?~; �/�?�/�?�?�?�?�? OO,ORO@OvOdO�O �O�O�O�O�O�O_*_ _N_<_r_`_�_�_�_ �_�_�_�_o&ooJo 8ono\o~o�o�o�o�o��o��EFPOS1� 1�̩  x�/:y�A?cN ��x-?y��� �"��F��C�|�� ��;�ď_�������� �B�-�f����%��� I��������,�ǟ P�b����I�����ί i�򯍯����L�� p����/���ʿe�w� �����6�ѿZ���~� �{ϴ�O���s��ϗ�  �2������z�eߞ� 9���]��߁����� @���d��߈��5�G� ���������*���N� ��K������C���g� ��������J5n 	�-�Q��� �4�Xj Q���q��/ �/T/�x//�/7/ �/�/m//�/??>? �/b?�/�?!?�?�?W? �?{?O�?(O:O�?�? !O�OmO�OAO�OeO�O��O�O$_�Cu2 1��O�O_�_{_�_ �O�_s_�_�_�_2o�_ Vo�_zoo�o9oKo]o �o�o�o�o@�od �oa�5�Y�} �����`�K��� ���C�̏g�ɏ��� &���J��n�	��-� g�ȟ��쟇����4� ϟ1�j����)���M� ֯q�����ϯ0��T� �x����7���ҿm� ����ϵ�>�ٿ��� 7Ϙσϼ�W���{�� ���:���^��ς�� ��A�S�eߟ� ���$� ��H���l��i��=� ��a���������� �h�S���'���K��� o���
��.��R�� v#5o��� ��<�9r �1�U�y�� �8/#/\/��//�/ ?/�/�/u/�/�/"?�/xF?,_>T3 1�I_ �/???�?�?�?�/O �?)O�?&O_O�?�OO �OBO�OfOxO�O�O%_ _I_�Om__�_,_�_ �_b_�_�_o�_3o�_ �_�_,o�oxo�oLo�o po�o�o�o/�oS�o w�6HZ�� ���=��a��^� ��2���V�ߏz���� ����]�H������ @�ɟd�Ɵ����#��� G��k���*�d�ů ��鯄����1�̯.� g����&���J�ӿn� ����̿-��Q��u� ϙ�4ϖ���j��ώ� ߲�;�������4ߕ� �߹�T���x����� 7���[������>� P�b������!���E� ��i��f���:���^� ����������e P�$�H�l� �+�O�sY?k44 1�v? 2 l��/2/�V/ �S/�/'/�/K/�/o/ �/�/�/�/�/R?=?v? ?�?5?�?Y?�?�?�? O�?<O�?`O�?OO YO�O�O�OyO_�O&_ �O#_\_�O�__�_?_ �_c_u_�_�_"ooFo �_joo�o)o�o�o_o �o�o�o0�o�o�o )�u�I�m� ��,��P��t�� ��3�E�W����ݏ� ��:�Տ^���[���/� ��S�ܟw� ������� ��Z�E�~����=�Ư a�ï���� ���D�߯ h���'�a�¿��� ��
ϥ�.�ɿ+�d��� ��#Ϭ�G���k�}Ϗ� ��*��N���r�ߖ� 1ߓ���g��ߋ��� 8�������1��}�� Q���u������4���X���|������5 1�M�_��� ;A�_���� �T�x�%� ��j�>� b���!/�E/� i//�/(/:/L/�/�/ �/?�//?�/S?�/P? �?$?�?H?�?l?�?�? �?�?�?OO:OsOO�O 2O�OVO�O�O�O_�O 9_�O]_�O
__V_�_ �_�_v_�_�_#o�_ o Yo�_}oo�o<o�o`o ro�o�o
C�og �&��\�� 	��-����&��� r���F�Ϗj�󏎏�� )�ďM��q����0� B�T����ڟ���7� ҟ[���X���,���P� ٯt�����������W� B�{����:�ÿ^��� ����ϸ�A�ܿe� � �$�^ϿϪ���~�� ��+���(�a��υ� ���D��߳���6 1���zߌ���D�/�h� nߌ�'��K����� 
���.���R������ K�������k����� ��N��r�1 �Ugy��8 �\��}�Q �u��"/��� /|/g/�/;/�/_/�/ �/�/?�/B?�/f?? �?%?7?I?�?�?�?O �?,O�?PO�?MO�O!O �OEO�OiO�O�O�O�O �OL_7_p__�_/_�_ S_�_�_�_o�_6o�_ Zo�_ooSo�o�o�o so�o�o �oV�o z�9�]o� ���@��d���� #�����Y��}���� *�ŏ׏�#���o��� C�̟g�🋟�&��� J��n�	���-�?�Q� ���ׯ���4�ϯX� �U���)���M�ֿq�x������7 1��� �����q�\ϕϛ��� T���x���߮�7��� [�����,�>�x��� ���ߘ�!��E���B� {���:���^���� �����A�,�e� ��� $���H�����~��� +��O����H� ��h��� K�o
�.�R dv�/�5/�Y/ �}//z/�/N/�/r/ �/�/?�/�/�/?y? d?�?8?�?\?�?�?�? O�??O�?cO�?�O"O 4OFO�O�O�O_�O)_ �OM_�OJ_�__�_B_ �_f_�_�_�_�_�_Io 4omoo�o,o�oPo�o �o�o�o3�oW�o P���p� ����S��w�� ��6���Z�l�~���� �=�؏a����� ��� ��V�ߟz����'���8 1�*�ԟ�  �����¯ȟ毁�
� ���@�ۯd�����#� ��G�Y�k�����*� ſN��r��oϨ�C� ��g��ϋ�߯����� �n�Yߒ�-߶�Q��� u�����4���X��� |��)�;�u������� �����B���?�x�� ��7���[�������� ��>)b���!� E��{�(� L��E��� e��/�/H/� l//�/+/�/O/a/s/ �/?�/2?�/V?�/z? ?w?�?K?�?o?�?�? O�?�?�?OvOaO�O 5O�OYO�O}O�O_�O <_�O`_�O�__1_C_ }_�_�_o�_&o�_Jo �_Go�oo�o?o�oco �o�o�o�o�oF1j �)�M������0��T�:�L�M�ASK 1�W��N�����x�XNO�  ������MO�TE  ǌ  ���_CFG ���O�l�PL_RGANG ��q[��A�OWER �W��y�`�SM_DRYPRG %W���%����TAR�T �q���UME_PRO������H�_EXEC_E_NB  �t\��GSPD��6�>��K�TDBY�k�R�Mz�k�IA_OP�TIONQ���^��INGVER-S��Ȋ
�o��I_AIRPUR�O� ��Մ1�m�M�T_��Tl��`�O�BOT_ISOLECŌ�-�4�0�o�/NAME���n��OB_CATEGňy�փ̀���س�ORD_NUM �?q�*�H769  �t�@�R�d�x�PC_T�IMEOUTQ� �xx�S232�1��ȅj� L�TEACH PENDAN���8����Ƽ ��pM�aintenance Cons�r�����"���tNo Use����π@�R�d�v߈�v���N�POΐ��8�̥ޙ�CH_L����^�J�	���!OUD1:1���R��VAIL!�¥�|\��SR  ��ʡ8���R_I�NTVAL����\��໮��V_DA�TA_GRP 2��ȅ�� D��PL�/�H�S�>�ȅ v���n����������� ������F4jX �|����� �0TBdfx ������// */P/>/t/b/�/�/�/ �/�/�/�/??:?(? ^?L?�?p?�?�?�?�? �? O�?$OO4O6OHO ~OlO�O�O�O�O�O�O��O __D_́�$S�AF_DO_PU�LS���p[��S'CAN}���[����SCm���`�Xj�+�p�p
��1�P`��վQ�r H� �_oo,o>oPo�_to��o�o�o�o�o�����ib2�d�Q�Qd�x�a
q�	�T�i @7�FXjtv&y�: ��t�_ @�sTʠ������T D���+�=�O�a�s��� ������͏ߏ����'�9�K��߯�8w�Z�����n�  =��;�o��ʑ��p����
�t��Di_�jaѰ�?X � ���� �U�Q9�K�]�o����� ����ɯۯ����#� 5�G�Y�k�}������� ſ׿�����1�C� U�g�yϋϝϯ���������	ߗ���2�D� V�h�zߌߞ߰���� �e�� ��$�6�H�Z�@l�~�����}�0�r ��&�������)� ;�M�_�q��������� ������%7I [m����� ��!3EWi {������� ////A/S/e/w/�� �/�/�/�/�/�/?? +?������ibk?}?�? �?�?�?�?�?�?OO 1O?IROdOvO�O�O�O �O�O�O�O__*_<_ N_`_r_�_�_�_�_�_��_�_oo&o8o,x� a��Co�o�o�o�o�o �o�o�o"4FX j|���zmo�\��v��+�����	12345�678]2h!B!��%�\1}�k`�T�f�x��� ������ҏ��lo� �1�C�U�g�y����� ����ӟ���	��-� >���a�s��������� ͯ߯���'�9�K� ]�o���@�R���ɿۿ ����#�5�G�Y�k� }Ϗϡϳ����ϖ��� ��1�C�U�g�yߋ� �߯���������	�� -���Q�c�u���� ����������)�;� M�_�q���B������ ����%7I[ m������� �!3EWi{ �������/ ///�S/e/w/�/�/ �/�/�/�/�/??+?@=?O?a?s?�?McE��?�?I/�?�?O�Cz  BpIj_   �H2_b� } �6F
[G�  	�AD�?�O�O�O�O�KDo�<�uO_$_ 6_H_Z_l_~_�_�_�_ �_�_�_�_o o2oDo Voho�O�o�o�o�o�o �o�o
.@Rd v�������D#��B�1iA�<�� �iA  �/�I��v,�mA>mAt  6@m�����x`�$SCR�_GRP 1��*P30� �� ��A ��	 Ё�؂�� �1����w��#��J��M�K@G�DC�v���N�G��L�	M-10iA/�8L 12345_67890k@��� 8k@MT20� ͐-C
ș�X��A^H �؁�Z�ǁ'�ǁ�C�G���-�	�v����������ά��H�؀_�܇ǂ���@�5�G���o�A"����������^� }h@,V�l\@-��B�%@��������A6@ �  @0�@8��N�?�^����H%@q�K��F@ F�`�£Ϛ��� ��������!��E�0� i����8�h�ߑ��ߵ�B���X�	��� -��Q�<�N��r�� ��������O�q�3�!�F��]@C�x��B<`�8�>���~�6��i�@8���%@����ȗ�'��?-DA!��1a�]�> �A	2�A T{��
�i���� (� � $��H3l)J��Γ��ECLVL  �A���7�?A���*SYSTEM*��@V9.1021�4 �8/21/{20�A �@��z�SERVE�NT_T   �$ $S_NA�ME !	 P�ORT�@!RO�TO! �_SP-D  ��/ �TRQ   �
,#AXIS5!�:'2  2c�,#D�ETAIL_ � l $DA�TETI! ER�R_COD�#IM�P_VEL4@ �	�"TOQ�$AN�GLES�$DIS���&" G%%$L�IN�" +$REC�5! ,!O%i � MRA�! 2w d2IDX�"��$B  �0$�OVER_LIM�I I 	 x,#O�CCUR5! � �+COUNT�ER�%FZN_C�FG5! 4 �$ENABL�#SyT� "FLAG"�DEBU�3R�! �V}4��5! �� 
$MIN_�OVRD�@$I��� �2�1�5FAC�Ee"�1SAF�7MIXEDL�9�!�2�ROB%$NE�&APP&4HELL��4	 5$�J?@BAS�#RS�R_�5  $�NUM_y@�  �xA1�'y@2�J3��J4�J5�J6�J7r�J8�'lAROO �� CO�ONLY��$USE_A�B#xBACKE�NB�  PIN>0T�_CHKSOP_�SEL_�0,Y_P�U;Qo1M_�!OU#PNS|F PYC�&��0EPM�%TPFWD_KAR�! P�!�RE$$OPT�ION�2$QUEԃY" D�RYRB$C�STOPI_AL;SYCEX+STQ�P�$[XTSPM1i2"�MA�1STY;TSmO
`NBRDIGQ�TRI�3�Q�WIN�I�M& 8bNRQ�xf`ENDNd$�KEYSWITCaH�S�QZa�THE�P�BEATM�SPE�RM_LE�"�QE�� �gU�SFd�RS~_dDO_HOM�09ORA/PEFP !"0L�3U ST�bRC�`�OM�#�!OV_M�SJQ ET_IOGCMN+S�W5aǀ�XEHK !
 D ��7qSU�"�RM�P+S� PO7B$�FORC�SWAR�NQ�XEOM�rP 7�$F'UNC��3U	0}QSAR'`�u2�v3�vY4�q��SC0O�P�L�r�"�XUNLiOeP�$:�ED� ���SNPX_�AS�2 0�@A�DD�0�1$SI}Z�!$VAR�'�MULTIPR�Z��pA�q �� $tY[�r	��B`�"�AC� ΆF'RIF">0S�P�y�"t��NF{dODBUS_ADw2�B���&CM�aDIA��q$DUMMY�15aM�3J�4J���Sz@  � Lx��"TEqM�8J��SGL��TAJp  &�0���@J�<����STMT�Q���PSEGb��BW<�P��SHOW��!�BAN̐TPOF��M�9J�0J�(a_��SVC�G�2; ��$PCpP?0\-�G3$FB�qPD�KSP�PAFPF�*��D/��2� ��!A0��@� �� �p���p��	������U5��6��7��8��9��A��B���p��h ��Ր��F���P����T�P���l�P�̩1�٩1�1�1 �1��1�1'�14�1BA�1N��!ǘ�2��U2��2��2̩2٩U2�2�2 �2�U2�2'�24�2A�U2N�3��3��3��U3��3��3̩3٩U3�3�3 �3�U3�3'�34�3A�U3N�4��4��4��U4��4��4̩4٩U4�4�4 �4�U4�4'�44�4A�U4N�5��5��5��U5��5��5̩5٩U5�5�5 �5�U5�5'�54�5A�U5N�6��6��6��U6��6��6̩6٩U6�6�6 �6�U6�6'�64�6A�U6N�7��7��7��U7��7��7̩7٩U7��7�7 �7�U7�7'�74�7A�Y7N�(2VP�`U3"� < �B
�*�� ! x �$TOR�Q@�  �"M$ R1 L@BQ_W0R��%T!�pJ�$S[C�Qp��_U���YSL|�   � x� ��7��m��0���`�R�VALU�5QP�V�]�F�ID_L��"%HI*I�r$FILE_xSM$BDk$s?�SA21� h5y E_BLCK�S�"���(D_CPU�)y��)�m��3P/b$��`sRR�  � PaWY0P�� 1LAƑ�S11314RUN_FLG(54,1�4�`/5M14M15H`rP4o04W�T2�Q�_LI�r  ]k@G_Ob�P�P_EDI+R��T2 @�3�20�$P��!����TBC2x� �}�8P/0T�Q�1FT'dD5cTDC/0A`a�0@aM	�F.AGTH�"��DDOPGRQH��pERVE(crD5c�rDa��0BC4PG@ X -$�ALEN(c�D5c�@`cRA�PF��W_k��#1�A:$2�GMO$�!C�S�DPIZP�`F!Y8�@![DE1U��LACEXrfCqCB���`_MA^�p0VjU@WjQTCVq\�Q@WT�a�Z�U�Zd��/S]��U@S]�J@`AG�M�T Jjgv�/U)a@U�A2)pp�\�5a.SH�JKHfV�K$�ZaU�Zaa�O`J��ra^cJJfcJJncAAL^c�`fc�`Ȏfm��b5OC�PN1��\�`�[nP�L
P_��� ��0CFb�{ `5GROU (���P�N�0C�� p?REQUIR]B��EBU̓�A�V$T1P2Vq�@@v�1�a��4 \�p�8A�PPRLpCL�
u$�0N�xCLO�0"�yS:E�y/U
�1�� ��0M,@oP�P�F��t_MGI��pC�x�z �d�lP�BR=K�NOLD��RTMO�1I�6��u	J�0H�P�dLPfcLP@ncLP�cLP�cLP6��97����V�2�5� Ir�B$���U��PATH ������H��p[p9�.�SCA�2L�l�r�qIN�BUCP��A\�Cf�UMe�Y�@k `l�&!xA�����������PAYL�OAD�J2LR'_AN$AȓL0ҙ�Αޑ�R_F2�LSHRlD�LO�Ӕ[��i��i�ACRL_�AY�L�U���r�bH��$H�^z�FLEX�s�1J�6 P�r�?
O�qO�O ���E  :�O�F@P�#���O�a@P�O�O�LF1 #�q����O__0_B_T_��E^_p_�_�_�_ �_�_�_�_�ȩ��Wc Hd����o!o3o"�:j	T�Ǌ�Xr��Fe�� �QeZ�3�]ooo�o�` �e�e�e�e�o�o�o�i8� ��t! ��00#5 AT��Hq��PEL�T1p�OxJ�[p VpJE3�CTRU���TN)l�@wHAND_VB�q�� ׄ" $���F2�<D�SW��b��0�v#� $$M��yM#���2�-�O� �q�K�A@) ���v(!h� �A��#�A1�A@�s��T� #�D1�D@�P �G"0		ST%�2�NC�DY.0�p� T�{����@�#���@��Hg��K�-�G�P�� ������������ʂ�bJ�5$ ����� Ʊ�qAS�YM0��Ip0�#wL��P�_n0A�a� t�^�`��~�������ƓJ͜~�ߚ����.��_VI��<(�sM V_UN�2; b#��
�JIez"�z"� ~$4��$�&=��PP�~�_�q�5;������Bf�0HR�0�1%��01���2DI@�;sOpO4ς10�& ��
��IeA��4�|1�����3��|��p�20 �' � ��M�E���Х2�"�TC0PT����1�`������8�1�9T���a $DU�MMY1��$P�S_��RF^��`u$(F�pFLAp�YP2�BB�3$GLB_T�E5]E�0ౡ�`۰��1( XX�p@wׁST��Vp�SBR�M21_�VRrT$SV_E�R�O��C�CCL�w@�BA�O2,0G�LD EWq) 4\p�1$Y��Z��!WS>`���A�0e�� 
�CU�E* ���N P�$G�I��}$�A p�@�CPq+ Lp\AV�}$F�EIV�NEAR�N��F��Y�TANC��C?�?�JOGR�t�� ,��$JO�INT=�N����AMwSETq-  >WEvU�:�SA�ZU;�q.� ��U���?�VpLOCK�_FO���K0BG�LV��GL:hTE�ST_XM�p�QEMP�PRr^buB%`�$U��B=�2*VpS�a+Ob��*`�a�)�ACE�`RS�` �$KARP�MQ3T�PDRA�@�d�QVcEC4��f�PIU�a�,�aHE,`TOOiLe��cVd�RE�`'IS3�r6�����ACH�P[p-qO�>��3D3��QPS�I�r  @$R�AIL_BOXEz=��@ROBOUd�?��AHOWWA�R��tq%@@qROLM0B�u �=t�r0�bp܍�ـO_F1�!>�@HTML5D1U�!0@�B2qځ/�^� R�`O��0�R]��Q��p!@��AOU�R1 d�@�e)�v�P�%`$PIPVfN 0�rbr2q���a�p�?CORDED*`6�L��PXTV�DQ),0�,�O�0 2 D \@OB��z�*`�����C[@���|�S;YS��ADR{�,0��0TCH:� 3� ,��EN52��A
1a_AT�	���+1�VWVA�14 Ǥ �`�BE5PR�EV_RT�$�EDITT�VSHWR1��Fs�� Q%< D�0�����?$HEAD�� 4���\�KE Q@�CPSPD��JM%P��LD5��R�g4�5�����I_`S{�C��NEp|��OTICKe�oM���`2�HN�A6 �@����Ñ_GP8R�Yv��STY	�>qLOwA,��0�N� �_7 t 
O�G�S%$4�AT=�@Sq�!$p!=м1HEy0rGFPRR�SQU�`xX�IB;!TERC�0���+0S�8  HP�@.�0�-���a^�1O�0�3��IZJDAQFE$APR��1Ap����.�PUAဵ_DYO�R�XS�PKD6�AXI���s�aURI��|�{p@�͆��J�_�`߂ET�P�3b��5(P�p6��A,B8D9Hw���$�)RSR��9l ��M�%�[�8�m� K�[�V�[�d�[�t��� ���Ŧ��Ŷ������������!��C6���C��ͯ����PTS�SC_@ : h��@DS`��a@SPLv0��AT��L����?��BADDRE�SsB_�SHIF�A�{`_2CH{�rɁI~@��TU~@�I*� ;�RCU�STO�*1VbI�j2< �Gh��d�
�^j
�rV-����0= \�@G����o�>��P��C��A��~�F���B���TXSCR�EE��><0��T�INA�COP��ATp%����? T�� �@d�߁�A�@L���ނ8��H�[�RRO �P`ހ��E�Ŵ��UE�G@ �-��6@S�AN߁RSM?���U��0
�D6��00S_S��@i������i�Cb���3� 2?��U�EAp2�Bp�G+MT� L�!���@�O�TC_�BBL�_BpW�0�0B �Ԟ�vOQ�LE��zpE�RIG�H�BRD�D�C'KGR�0�T���>�WIDTHHs���Ĳ!ABAq�UMI�pEY�Щ1C6���p�p��bpl�BACCK��0B1�A�0sFO�DLAB���?(�0I@p#b$�UR�qq�
�0H>l� D 81�P!_����0R P%b /�Hx Aa0�O�0%EI��G� U� �9R3b�qLUM�Ķ��ERVM�N�
PԔPF�0�GE`u{Q������LP4%
�E���)Q'��_(P��_(,p^)5\+6\+7\+8A"��3k��P���F,qaS�P�E	USR�DG <�@�0UERT�ERsFOB�ERPRI��mLp�!30TRIP�^qm�UNDO
g5H<PàL0���qƤ��{bްؠ qI�� o�G ��aT�p�� �2OS�1��6R�r�v3�a�AJ��OS^�2b��P{bU<!�AK�?�?��<"a�Nv3OFFT`�@L�@��3OU@ 1Jh�@?DgDK�@GUف�PfA�R�C}ьGS�UBb��@/ SRT��0B�MI��Q�pO�O9RBp�ERAUT��D�T�I��A_R��Ns |]��OWNy0>�$SRC}������DT`>UR�MPFqIy�y��ESP|��G��u#��'r��Um�6O `@W�O���=��COMP!A$հ{0_YP�r�Q.��UWA_�C ra�Q�P�S�Qr��4�ܘrW� P?�SH�ADOW��s"a_UNSCA�c"c��/cDGD7q��EG�AC�Sd狠PPG��Q���STEĉ��O��t�PEZ"��VWDt}�TRG�6R �<>��jMOVE}����bANG���f-C�f|�3�bLIM_X!C v'Cv�hq|��g0?06��`��VF���CN�VCC���S?�C��RA���`ϥD�.�@NFA�R@�]�-E,�Q>0G����R:�{0DE�b��p���p6T� i�؁ϣ�u���W C% �DRI�`��aV[�*��S��D�$MY_UBY �$�}�3ϥ~���1��a��P_8`y�ڶ�L��BM�$n�DEY
�EXc ,���UMUِX�d�����US��˰.0_R����#06��fG�PACIqt�`HQ�dI��-CI��3I����QRE���1�B�sI�U ?�PG�`P��⎐t0�sR�0�V �k���B	�R���R�dSWA�os�@$��n�O�!�A���[�E� U���a�@��0�sHK��W����aS���Q��cEA�NS��P�����rMwRCV6X �- UO�pM�C��	��8?C����REFb�� ����
r�ِ0���@��꡹����A�_;P W�B�o����`��k�\����x��A�r3Y ���a��ϒ�1`�$GROU���3��¶��s�pT����20$0 ����0X V�Ӂ�Xֱ���UL�qW�P�C%p�X��NT�S+�b*��6��!6���L��_Ű�_���k��!�pTIЙ�Z� t@MD�@AP�_HUx��`��SA.�cCMP}�F�����Ų�_��Rqty����W�j�X�ɗQVGF|`S[� �qM0����UF_{�0˂��@JʼRO� T��շ����|.�UR1E9��6�RI;���I&༨�o�o{FQyXFQ'C`wIN�H��xx� V�1,r��A��?�W�|��Q/��V����LOp'�\ax ������!NSI"V�IA_�R;�\ ��� HDR )�$JO� b��$Z_UP)p��Z_LOW�������\(p���P鱬3�9���Ⴐ��'Q��p| �"�]� 0��PA� �CACH���}���퀙��!�P]SC(qIB�F�#���T� ��|�$H	O�1R��/�%�" f������?�RQ0!���cPVP��� H_SIZ�RZ��M��N�Q�MPr
�qIkMG�d��AD�	��RMRE���WG�PM�pNDRP�VA�SYNBUF�VV�RTD� W��OLE_2D,tc�J1@C�qUۃ��Q���ECCU{�VE�Me�}�d��VIR�C��
" {�L�A��RQ}0\0��AG:R�XYZ)��C�W�������A�T�p܂IM��|G`��GRABB�1�Y�b�� ���^�>
�CKLAS��8b�Y@_  񱵵IT��5P@�21T$b��p!�` ���SP�G�%TQ�RQ�q�P�"�x�I�$|��=�BG�_LEVE�QL�PaKL��"ѥ�GI� �NO�Q܁��"H�ObPRa �  �F����E6S��g�]2RO�cACCE0e@����x4VR�A`�y1܂R`� AR�c�PA@�>��D�SRoEM_BQ$ ��N͐JMPU�XAbi$�1�$SSlSO�
���S�G�Y@c � ��S� ��N\/D��LEX�&db`Sdqg`��&DR�w�$YQqH(`qH҄�cޞ��VP2h�e'� �є`V��cPMV_PI��DX �`�@3����IF&�\rZ�JT�E�@���H����E�AGAU?�LO9O�d?�JCBTZ�'�B`H +cPLAN'r��L2��Fw��D?V5Y �WM��~Ppu�T�FS��U�Q�ѥU@����V2DbX�1�LRKEZq�1VAsNC]C`�R_O�|`f (�p8�s$p\�3Zr�rR_A3� g 4��dovn�#p� çB��h h���9��ĬvOFF��sfW@�����EA���
� LSK��M8N��q�g S`��||@c"i < WJ���=�UMMYY�j��n�D�Pȉ!�CU��1�U�pj� $�TITV1�$PR8A��OPL����SF���Cki ��|6���)1SMEO!�l%BXC�4J�p���ZD�vm DlQx�AL^1IM; ���0IN�MSG_Q�Sw@�I_pn%B�w8�x%�M� �XVR"��oI"�pT�5���ZABC��p�Ƃ��Ӡ
)��%��`VS.� q � w0���=�CTIVeAI�O�b�	s�ITVlLW�DV@
l�"��2� DI�� @�� ��|A��d���N�LSTs���ݰ���_ST��	C}_�DCSCH��r LQp�����~P01��m�W GN����xr���_FUN��� A04�ZIP�!�s%B� L8�L�|�Ѣ�AZMPCFʅt�r9���L�?DMY_LN$pq�7�'�˄u �$��Q�CMCM���CLCART_���P�a $J����D=��¢ ��u�ǥu���_�p����UX�P�UXEUL����
��̥
��.��>���FTF���k���7��Cv_��*�����Y%�D.  w _8 $R� U�Q���EIGHe3�x?(�0��0�� ��A$�x �=0�s���$�B�����b_SgHIFB�	�RV�P�F��1�	$)0C �ঢ���d�pl��rH�"l��D|ȕ�C ��NV�a��SPH�0%�y ,�0��ֿ���$S{0DE�FAUn��b����_�����'HOT�������MIPOWERFSL �B����%�oWFDO�� ��� ��Y��`1 ����q�� L!=ip_EIP5ԑ�~���j!AF��x�`�߼�!FT��2�����!��-�s���S�!R9MHQp�7�B��f��@o�5黎���!�OPCUA���y��7�!TPPȜ@8���d&���!
3PM�p�pXY����Aer���J����f���!RDM-@V���g
g!R�90h��hV�!!
h�~�����i���!RLSYNC� &8�K!gROS��r�4:ޗ!
CEL�MT��`���k��!	$��PS���l�//�!�WASRCd6��m/{/!�'USB|/��nj/�/!STMP��/��o�/?�7?*?`=�e�I��KL ?%�q� (%SVCPRG1`?�:�52�?�?�03�?�?�04�?�?�05 O%O�06HOMO�07pOuO�0�8�O�O�09�O�K �4~�O�1�?_�1�? =_�1�?e_�1O�_�1 :O�_�1bO�_�1�Oo �1�O-o�1�OUo�1_ }o�1+_�o�1S_�o�1 {_�o�1�_�1�_E �1�_m�1o��1Co ��1ko��1�oe?w2 �0~?�00�u��1y��� �������Џ	��-� ?�*�c�N���r����� ϟ�����)��M� 8�q�\�������˯�� �گ���7�"�I�m� X���|�����ٿĿ�� ���3��W�B�{�fπ�ϊϱ�������k:_�DEV q���MC:�4����GRP 2�q����0bx 	� 
 ,c��|�<�hߥߌ��� ��������#�
�G�Y� @�}�d������� ���d�1���U�g�N� ��r�����������	 ��?&cJ�� ������� ;M4qX��� ���/�%//I/ 0/B//��/�/�/�/ �/�/�/�/3??W?>? {?�?t?�?�?�?�?�? O�?/OAO�/eOO�O �O�O�O�O�O�O�O_  _=_$_6_s_Z_�_~_ �_�_�_�_HO�_'o�_ Ko2ooo�oho�o�o�o �o�o�o�o#5Y @}dv�
o�� ���1��*�g�N� ��r��������̏	� ��?�&�c�u���� P���ϟ���ڟ�)� �M�4�q�X�j����� ˯�����%�|�� [���f�������ٿ �������3��W�i� Pύ�tϱϘϪ���7�d ���	���	��B�-�f�Qߊߙ�%�x�߾�>������ ������������9� '�]�k�ߐ���S�� �����������;�}� b���+����������� ����C�i�:y�m [����  ?�3�CiW� {����/� ///?/e/S/�/��/ �y/�/�/?�/+?? ;?a?�/�?�/Q?�?�? �?�?O�?'Oi?NO`O O9OO�O�O�O�O�O �OAO&_eO�OY_G_i_ k_}_�_�_�__�_=_ �_1ooUoCoeogoyo �o�_�oo�o	�o- Q?a�o�o��o �����)��M� �t��=���9���ݏ ˏ��%�g�L���� �m�������ٟǟ�� ?�$�c��W�E�{�i� ������կ���;�ů /��S�A�w�e���ݯ ¿Կ��������+�� O�=�sϵ���ٿc��� ��������'��Kߍ� r߱�;ߥߓ��߷��� ����#�e�J���}� k��������+�Q� "�a���U�C�y�g��� �������'����� +Q?uc���� �����'M ;q���a�� ��//#/I/�p/ �9/�/�/�/�/�/�/ ?Q/6?H?�/!?�/i? �?�?�?�?�?)?OM? �?AO/OQOSOeO�O�O �OO�O%O�O__=_ +_M_O_a_�_�O�_�O �_�_�_oo9o'oIo �_�_�o�_oo�o�o�o �o�o5wo\�o% �!������ O4�s�g�U���y� �������'��K�Տ ?�-�c�Q���u����� ���#�����;�)� _�M���ş����s��� o�ݯ��7�%�[��� ����K�����ſǿٿ ���3�u�Zϙ�#ύ� {ϱϟ��������M� 2�q���e�S߉�w߭� �߽��9�
�I���=� +�a�O��s������ ������9�'�]� K��������q����� ����5#Y��� ��I������ 1sX�!�y �����9/0/ �	/�Q/�/u/�/�/ �//�/5/�/)??9? ;?M?�?q?�?�/�?? �?O�?%OO5O7OIO O�?�O�?oO�O�O�O �O!__1_�O�O~_�O W_�_�_�_�_�_�_o __Do�_owo	o�o�o �o�o�o�o7o[o�o O=sa���� �3�'��K�9� o�]�����̏��� ���#��G�5�k��� ����[�}�W�ş��� ��C���j���3��� ������������]� B����u�c������� �����5��Y��M� ;�q�_ϕσϥ���!� ��1���%��I�7�m� [ߑ��ϸ��ρ���}� ��!��E�3�i�ߐ� ��Y����������� �A���h���1����� ����������[�@ �	sa���� �!���9 o]����� �/�!/#/5/k/Y/ �/��/�/�/�/? �/??1?g?�/�?�/ W?�?�?�?�?	O�?O o?�?fO�??O�O�O�O �O�O�O_GO,_kO�O __�Oo_�_�_�_�_�_ _oC_�_7o%o[oIo ko�oo�o�_�oo�o �o3!WEg� �o��o}���� /��S��z���C�e� ?����я���+�m� R������s������� ߟ͟�E�*�i��]� K���o�������ۯ� �A�˯5�#�Y�G�}� k����	�ڿ���� ��1��U�C�yϻ��� ߿i���e���	���-� �Qߓ�x߷�A߫ߙ� �߽������)�k�P� ����q������ ���C�(�g���[�I� �m�������	���  ������!WE{i �������	 SAw��� g����/// O/�v/�?/�/�/�/ �/�/�/?W/}/N?�/ '?�?o?�?�?�?�?�? /?OS?�?GO�?WO}O kO�O�O�OO�O+O�O __C_1_S_y_g_�_ �O�__�_�_�_o	o ?o-oOouo�_�o�_eo �o�o�o�o;}o bt+M'��� ���U:�y�m� [�}����Ǐ���-� �Q�ۏE�3�i�W�y� {���ß��)���� �A�/�e�S�u�˟� ¯��������=� +�a�����ǯQ���M� ˿�߿��9�{�`� ��)ϓρϷϥ����� ���S�8�w��k�Y� ��}߳ߡ�����+�� O���C�1�g�U��y� ������������	� ?�-�c�Q������������$SERV_MAIL  ��������OUTP�UT�����@��RV 2vw�  �� (�x��I��SAVE���TOP10 2}#	 d �� �����' 9K]o���� ����/#/5/G/ Y/k/}/�/�/�/�/�/ �/�/??1?C?U?g?`y?�?�?w�{YPf���FZN_CFGw w����W�1GRP �2�7t ,B�   A'@��D;� B(@�  �B4�RB2�1VHELL�2!	w�r6 7�7�O>�K%RSR�O�O �O�O�O_�O3__W_ B_T_�_x_�_�_�_�_��_on�  ���RoKo]o+bio ���eo�b�`�bg3b2��dultm�b�RFHK 1
`K �o0Y Tfx����� ���1�,�>�P�LL?OMM `O���QBFTOV_EN�B��+r�bOW_?REG_UI�����IMIOFWDL⋀��*E��WAIT���i�2���ᆹ*�TIM���T�VA��+���_UNIT����r	�LCڀTRY��r��MON_ALIAS ?e��2 he���!�3� E�S���v�������W� Я�����ï<�N� `�r���/�����̿޿ 𿛿�&�8�J���[� �ϒϤ϶�a������� �"���F�X�j�|ߎ� 9߲��������ߥ�� 0�B�T���x���� ��k�������,��� P�b�t�����C����� ������(:L^ 	�����u�  $6�Zl~ ��M�����  /2/D/V/h//�/�/ �/�/�//�/
??.? @?�/d?v?�?�?E?�? �?�?�?O�?*O<ONO `OrOO�O�O�O�O�O �O__&_8_J_�On_ �_�_�_O_�_�_�_�_ o�_4oFoXojo|o'o �o�o�o�o�o�o 0B�oSx��� Y������>� P�b�t���1�����Ώ ��򏝏�(�:�L��� p���������c�ܟ�� ��$�Γ�$SM�ON_DEFPR�OG &����N� &�*SYSTEM�*+�o�����?=�RECALL� ?}N� ( ��}!xyzra�te 124=>�169.254.���120:19636 ��ɠȡ���l��}
��1 �� ǯٯj�|���!���;� ��_����'�ο˿ ݿnπϒϥ�L�I�[� �����#ϵ�����j� |ߎߡϳ�E�W����� ��1�����f�x�� �߯�A�S������� -������t������ =���a�����)��� 8��p����NK ]� %��� l~��5GY� �/!3��h/z/ �/��C/U/�/�/
? ///�/�/d?v?�?�/��/??Q?c?�?O=:�copy frs�:orderfi�l.dat vi�rt:\tmpback\�?�2dOvO�O;1*Bmdb:g*.*?OQO6 \O��O�O_$25x*D:\�O4P�O�2�Oq_�_�_}6*Ua2_D_�? �_�_oO1O�OUOfo xo�o�O�OJo�O�o�o _-_�_Q_�ot� �_�_<Na����8 ���k�}�����?�?17572 �?]�� ��%?��ɏ�ۏl�~���#imd:�picksim_�part1.tp�eemp�oF���� �����?�̟ޟo��������tpdisc 0N�G�I�[��������tpconn 0 ϯůׯ�h�z�����2��omay��P�I�]�� �ϥ�2��ɿۿl�~���#�d��E�W����� ߟϱ�6�����k�}� ��"o4o�oX������ �o�o��F���m�������$SNPX_�ASG 2�������o  0��%������  ?���PA�RAM ����� �	��Pʠ�����1������OFT_K�B_CFG  ������OPIN_�SIM  ���,����������R�VNORDY_DOO  6�b����QSTP_DSB�v�,���SR ��� � &�0�Q����G�TO�P_ON_ERR�����|PTN ���� �A��RING_PR�M���VCNT_OGP 2x�.���x 	
	���0�T��VD� RP' 1�/�E�� 7������� //1/C/U/g/y/�/ �/�/�/�/�/�/	?? -???Q?c?�?�?�?�? �?�?�?�?OO)OPO MO_OqO�O�O�O�O�O �O�O__%_7_I_[_ m__�_�_�_�_�_�_ �_o!o3oEoWoio{o �o�o�o�o�o�o�o /Ahew�� ������.�+� =�O�a�s��������� ͏����'�9�K� ]�o���������ɟ۟ ����#�5�G�Y��� }�������ůׯ��� ��F�C�U�g�y��� ������ӿ��	���-�?�Q�c�mPRG�_COUNTW�9���ENB����M��Y���_UPD� 14T  
xϣ���/�X�S� e�wߠߛ߭߿����� ���0�+�=�O�x�s� ������������ �'�P�K�]�o����� ������������(# 5Gpk}��� �� �HC Ug������ �� //-/?/h/c/ u/�/�/�/�/�/�/�/ ??@?;?M?_?�?�? �?�?�?�?�?�?OO %O7O`O[OmOO�O�O��O��_INFO {1����P	 �O__@_�+Y@l�@Iʟl?Z�F_-S��̵��5A�u�9	�]�Ǝ�@�K]�A���@CP A!" ?�nn_��A D5Oy����C����($6�T�5+���Q� �8�h�Ca���.~:��1�５���YS�DEBUG�������@d��
`SP_PwASS��B?k�LOG �F.�  �@�X�O�  ����AU�D1:\Hd�NIb_MPCNm���o�o����a�o ���fSAV Qi��2Qqal�b�E�hSV�k�TEM_TIME� 1Qg� 0o`2T��Z����^sMEMBK  	����q`qo��� �X|��� @ ��C�"�G�W���z�����a 2[@}q��я���/s���1�C�U�g�y� �{�����ß՟�����/�i�e>�c�u� ��������ϯ��� �)�;�M�_�q���������\uSK�p�x��`������.�@e���2,�W�AW�A�����i��Ϧ�(��#!������� ���<�-�� �-���0`F�t߆ߘߌ�Y΀��������(��@$,�P�D�t��� �����������(� :�L�^�p��������������T1SVGU�NSPD2e '�e���2MODE?_LIM �vvqd b��2��Qm���ASK_OPTGION`�y aS�_DI+`ENB � b�esBC2_GRP 2ܵ c|r�[R��C������BCCFG �7| (��b�L_U@R� v������/ -//Q/</u/`/�/�/ �/�/�/�/�/??;? &?_?J?�?�?7ց<�? �?�?�?p?�?+OOOO :OsO~�O�th@�O�O �O�O�O	_�O-__=_ ?_Q_�_u_�_�_�_�_ �_�_o)ooMo;oqo _o�o�o�o�o�o�o�h �03EW�o{ i������� ��A�/�e�S�u�w� �������я���+� �;�a�O���s����� ͟��ݟߟ�'��K� c�u�������5�ۯ ɯ����5�G�Y�'� }�k�����ſ��տ׿ ���C�1�g�Uϋ� yϛ��ϯ�����	��� -��=�?�Q߇�u߫� a����������;� )�K�q�_����� �������%��5�7� I��m����������� ����!E3iW �{����� ��#5Sew�� �����//� =/+/a/O/�/s/�/�/ �/�/�/?�/'??K? 9?[?�?o?�?�?�?�? �?�?�?�?OGO5OkO !�O�O�O�O�OUO�O �O_1__U_g_y_G_ �_�_�_�_�_�_�_�_ 	o?o-ocoQo�ouo�o �o�o�o�o�o) M;]_q��� �O���%�7��[� I�k������Ǐُ�� ���!��E�3�U�W� i�����ß���՟� ���A�/�e�S���w� ��������ѯ���+� �C�U�s�����������˿�߿���3���$TBCSG_G�RP 2���  �3�� 
 ?�   ^�p�Zϔ�~ϸϢϴ�@�����$�7�>�E̿d0 �S�?�3�	 HCA��"�>l�"�CS�BpVߙ�c�u߇����B�$�>������"�Bl����)�A������G�"�;�B�)�+�Q�G��$_��A3�"�Q���T��Ѩ��@����� '�:���e���M�_�x������?�ff��� ��	V3.0}0V�	mt2 * 2�$��<23�G�� [ -\  q��7�+J2>�E����CFG !��eO� R��
����0� 0Vd�d�u� �����/// P/;/t/_/�/�/�/�/ �/�/�/??:?%?^? I?�?m??�?�?�?�?  OOV�p�O/OAO�? tO_O�O�O�O�O�O�O �O_(_:_L__p_[_ �__�_�_3���_�� �_ooIo7omo[o�o o�o�o�o�o�o�o 3!WEgi{� �������-� S�A�w�e�����m�ŏ ׏������=�+�a� O���s�����͟ߟ�� ���9�'�]�o��� ��M�����ۯɯ�� ��5�#�Y�G�}�k��� ����׿ſ����� C�1�S�U�gϝϋ��� ������	����?�� W�i�{�%߫ߙ߻߽� �����)��M�_�q� ��A��������� �%���5�[�I��m� ��������������! E3iW�{� �����/ ?AS�w��� ����/��O/=/ s/a/�/�/�/�/�/�/ ??�/%?K?9?o?]? �?�?�?�?�?�?�?O �?!OGO5OkOYO�O}O �O�O�O�O�O_�O1_ _U_C_y_g_�_�_�_ �_�_�_�_o	o+o-o ?ouo��o�o�o[o�o �o�o;)_M ����w��� ��7�I�[��'��� �����ُǏ���� 3�!�W�E�{�i����� ����ß�����A� /�e�S�u��������� �ѯ���o1�C��o ����s�����Ϳ��ݿ ��'�9�K�	�ρ� oϥϓ��������Ϲ� #��3�5�G�}�kߡ� ���߳��������� C�1�g�U��y��� ������	���-��Q� ?�a���u���%�W��� ������M;q _������� #%7m� �]����/� /!/3/i/W/�/{/�/ �/�/�/�/?�//?? S?A?w?e?�?�?�?�? �?�?�?OO=OOO�� gOyO�O5O�O�O�O�O �O�O_9_'_]_o_�_ �_Q_�_�_�_�_�_�^�  %`)c �)f=o)b�$TBJ�OP_GRP 2�"�U� _ ?�)f	Ub�\c$cl��P��pJ�`��xe  � �� � ��`�)d� @%`tb	 ��CA��f��S�C��_)eta�b3�33�f�oz=�_��CS�?��Y�1ru`B�;pp�gLWw�o�o?�a�u�ޜz<؄-r��a��u=�)eB��w?C�  D�a�o�#�-�;��B9l�`2u�ff�n�&)eAЇ��w���>��ͭ�����;�ǎ���@fff���b�]���A���������9�ˌ�X��@�o�폎������%��ɟۛ;������@�o��� {����9�1�g�Y�C� Q������E�ϯ�ӯ ��@��կ_�y�c�Pq���пct�)f���	V3.00�zcmt2��*��yd$a)�4� �F� G9| �G�v�G�/��G�� H�@�H,�H.���HC� HYA@�Hn��H�� �H�� H�Y@�H�`H����H�c�H��H̿�H�nD��G G.A �GKm Gh� �G��G�x��G��G����G�:�G�Ѐ�G�f�G����G��\��H
�_�H��H���H @�H'��d�ր=L��=#�
������)bQ3o�+�)f/��?�߀f�d�RcESTPARS�hn`�RcHR��ABLEW 1%ci�)d�_�D� �@$�_�B_�_�(g0a_�	_�E
_�_ؾ�)a_��_�_�����RD	I��ma�����������O������������S��kc  I���������� *<N`r��� ����Hm���� lb��C,�>�P�b�� �2�D�V�h��)N�UM  �U*ma�`1` ������_CFG &�+��a@U`IMEBF_TT�Ѻkc��T&VER�Uj&�T#R 1'��' 8&�)b$`�! �PN  �/�/�/ �/�/	??-???Q?c? u?�?�?�?�?�?�?�? <OO)OrOMO_OuO�O �O�O�O�O�O�O__ %_7_I_[_m__�_�_ �_�_�_�_4oo!ojo EoWomo{o�o�o�o�o�җ!_!�&@�%���MI_CHAN�`' �% .sDBGLVL`'�%��1p�ETHERAD �?���p�/���o�o��y�1pRO�UT~ !�!��t��|SNMAS�Kyx�#�q255.?��=�O�a�Á��OOLOFS_D�I���ecyORQCTRL (�+��0�ߍTΏ��'� 9�K�]�o��������� ɟ۟����#�3�͏�V�E�z�~�PE_D�ETAIWx��PG�L_CONFIG� .)"!���/cell/$C�ID$/grp1�~�����*�<��� �g�y���������P� ���	��-�?�οc� uχϙϫϽ�L�^��� ��)�;�M���q߃� �ߧ߹���Z����� %�7�I��������������M}n��!� 3�E�W�i��k���p��m���������  g�DVhz��- ����
.� Rdv���;� ��//*/�N/`/ r/�/�/�/�/I/�/�/ ??&?8?�/\?n?�? �?�?�?E?�?�?�?O "O4OFO�?jO|O�O�O �O�OSO�O�O__0_ B_�Of_x_�_�_�_�_��_͠�User View ��}}1234567890oo'o9o�Ko]oed�`£�o���Y2�Yb_�o�o�o�o !�o�o�R3�oo �����(��n4^#�5�G�Y�k�}�����n5�׏���@��1���R��n6Ə ��������ӟ�D���n7z�?�Q�c�u����������n8.�����)�;�M���n�t� �lCamera�Z꯳�ſ׿������E��7�I� [�ouχϙϫϽ���ŉ  ���i���1� C�U�g�y� ϝ߯��� �����	��-�?�f����]y�ߋ����� �����	��-�x�Q� c�u�������R�d�� B���	-?Q�� u�������� ��d��˰ew ����f��/ R+/=/O/a/s/�/, ��y�/�/�/�/?? )?�M?_?q?�/�?�? �?�?�?�?�/d�-��? ;OMO_OqO�O�O<?�O �O�O(O__%_7_I_ [_Od���O�_�_�_ �_�_o�O%o7oIo�_ moo�o�o�o�on_�W9So,>Pb 	os��Qo������(�:�ɪ	��0 �u���������Ϗv ����;�M�_�q� ����<�N�����9��  ��$�6�H��l�~� ��۟��Ưد���� ����ۥ�Z�l�~��� ����[�ؿ���G� � 2�D�V�h�z�!�[�n� ���������� �ǿ D�V�h߳όߞ߰��� ���ߍϟ���}�2�D� V�h�z��3߰����� ���
��.�@�R��� ��F����������� ����.@��dv ����e��Ų+U 
.@Rd� ������//<*/�  �	Y/ k/}/�/�/�/�/�/�/x�/?;   // 7/U?g?y?�?�?�?�? �?�?�?	OO-O?OQO cOuO�O�O�O�O�O�O �O__)_;_M___q_ �_�_�_�_�_�_�_o o%o7oIo[omoo�o�#<  
� (  ��M ( 	  �o�o�o�o�oC 1SUg����t��j?: �y *�<�N��r������� ��̏������a� >�P�b�t�����ߏ�� Ο��'���(�:�L� ^����������ʯܯ � ��$�k�}�Z�l� ~�ů����ƿؿ��� C� �2�Dϋ�h�zό� �ϰ���	�����
�Q� .�@�R�d�v߈����� ������)���*�<� N�`�߄������� ������&�m�J�\� n�������������� 3�E�"4F��j| ������ S0BTfx�� ����//,/ >/P/���/�/�/� �/�/�/??(?o/L? ^?p?�/�?�?�?�?�? �?5?O$O6O}?ZOlO�~O�O�O�O�?�p@ A�B�O�O_�C�G��`��#frh:�\tpgl\ro�bots\m10�iaAS_8l.xml�Oe_w_�_�_�_��_�_�_�_on�� o>oPoboto�o�o�o �o�o�o�oo: L^p����� �� ��6�H�Z� l�~�������Ə؏� ����2�D�V�h�z� ������ԟ���� 	�.�@�R�d�v����� ����Я�����*� <�N�`�r��������� ̿޿���&�8�J� \�nπϒϤ϶���������� XVA |�O+P<< )P ?���A���9�[� ��oߑ߿ߥ������� ���=�#�E�s�Y������������6��$TPGL_OUTPUT 1	A�	A !� -�B�T�f�x������� ��������,> Pbt�������-�!Є��2345678901 );M_g�2 ��������@/0/B/T/f/�}p/ �/�/�/�/�/x/�/? (?:?L?^?p??~?�? �?�?�?�?�?�?$O6O HOZOlOOO�O�O�O �O�O�O�O
_2_D_V_ h_z__�_�_�_�_�_ �_�_�_.o@oRodovo �o o�o�o�o�o�o �o<N`r� .������� "�J�\�n�����*����ȏڏ�������} �F�X�j�|��������@#�՟�)� ( 	 ��
�@� .�d�R���v������� �Я���*��N�<� ^���r�����̿��� ޿ ���J�8�n����8�vϨϺ͒��� �����$��
��U�g� �sߝ�w߉�����C� �����Q�c�=�� ���߁���i���� ��;�M���5�����/� ��������_�q�7 I��QYk�� %����3 i{���K�� ��///�/e/w/ /�/�/�/�/�/A/�/ ?+?�/O?a?;?M?�? �/?�?�?y?�?O�? OKO]O�?aO�O-OO �O�O�O�O_oO�OG_ �O3_}_�_i_�_�_#_ �_�_o�_1oCooOo yo�_�_�o�o[o�o�o �o�o-?�ocu�a�������)�WGL1.XM�L��(��$TPOFF_LIM ��|�����6��N_SV>�  ���P�P_MON7 2��R������22�STRT?CHK 3��P��C�9�VTCOM�PATe��T�VW�VAR 4��\�i� Ə *��I���:�_DE�FPROG %���%PART1 TLd�{���4��_DISPLAY�E���Z�INST_�MSK  �� ���INUSER�叜�LCK�QUICKMEN�ޜ�SCRE1������tpsc@���L�Q�P�b�_f��ST�P�RACE_CFG 5����I�	3�
?����HNL 26i�b�ѡ� ?��� )�;�M�_�q�������ITEM 27�� �%$1234567890ؿ�  =<���"�  !(�0�<��u�3�ֿ������ ��0���T�f�/ߊ�J� ��Z߀������4� >߸�b��4�F��j� ������l�������� ^������*�x��� �������6�H�l� ,��Pb��x��< � �D�(� 4���N��� �@ /dv�/$/ �~/�/��//*/�/ N/?r/2?D?�/Z?�/ �/�??�?&?�?�?~? n?�?�?�?�?0O�?�O �O�O"O�OFOXOjO�O �O:_`_r_�O~_�O_ _�_�_T_o&o�_2o �_�_�o�_�oo�o�o >o�obo�o=�oX�o h���(:L �p�B�T��x�� � �����6����l� �����k�Ə��ꏪ���� �ҟD�V����S�8��$��  ��$� ɡ{�r�
 ������үS��UD1:\߬���6�R_GRP �19Ż� 	 @{�*�<�&�\� J���n��������˿�ٺ��߯��'��?�  B�T�>�t�b� �φϼϪ�������� �:�(�^�L߂�pߒ߆��	�����4�S�CB 2:@� -�*�<�N�`�r������*�UTOR?IAL ;@�Ư��/�V_CONFIG <@�ġx��¯d��OUTPU�T =@�U���p�����������  2DVhz� R�������  2DVhz�� �����
//./ @/R/d/v/�/��/�/ �/�/�/??*?<?N? `?r?�?�?�/�?�?�? �?OO&O8OJO\OnO �O�O�?�O�O�O�O�O _"_4_F_X_j_|_�_ �O�_�_�_�_�_oo 0oBoTofoxo�o�o�_ �o�o�o�o,> Pbt���o�� ����(�:�L�^� p��������ʏ܏�  ��$�6�H�Z�l�~� ����>�P������� �(�:�L�^�p����� ������ܯ� ��$� 6�H�Z�l�~������� ůؿ���� �2�D� V�h�zόϞϰ���ӿ ����
��.�@�R�d� v߈ߚ߬߾������� ��*�<�N�`�r�� ������������ &�8�J�\�n������� ����������"4 FXj|���� ����0BT fx������ �//,/>/P/b/t/ �/�/�/�/�/��/? ?(?:?L?^?p?�?�?�?�?�?������?�?�1�?&OɟJO \OnO�O�O�O�O�O�O �O�O_"_�/F_X_j_ |_�_�_�_�_�_�_�_ oo0oA_Tofoxo�o �o�o�o�o�o�o ,=oPbt��� ������(�9 L�^�p���������ʏ ܏� ��$�6�G�Z� l�~�������Ɵ؟� ��� �2�C�V�h�z� ������¯ԯ���
� �.�?�R�d�v����� ����п�����*� <�M�`�rτϖϨϺ� ��������&�8�I� \�n߀ߒߤ߶�����������"�4�C��$�TX_SCREE�N 1>�5;�0�}�C�� ��������u�2F t�!�3�E�W�i�{��� ������������� /��Sew��� $�H�+= O������� �V/z'/9/K/]/ o/�/��//�/�/�/ �/?#?�/�/Y?k?}? �?�?�?*?�?N?�?O�O1OCOUO�?yO�$�UALRM_MS�G ?c��p� qOFګO�O�O�O_ _6_)_;_Y___�_�_�_�_�_�ESEV � �M
f�BE�CFG @c��m�  F�@��  A:a   B�F�
 �_M�c� moo�o�o�o�o�o�o��o!/waGRPw 2A k 0F��	 Woy�@I_�BBL_NOTE� B jT���lM�h�O��,`�rDEFPRO��@%�K (%�PART2z�|% �_��?�*�c�N��� r��������̏��{�FKEYDATA� 1Cc�cpp 	/gF�fi�{�R�������,(���F�(POINT�z� ҐIREC��B�)�ND-�l�'�C?HOICE]p���TOUCHUP ����ȯ�ӯ���4� F�-�j�Q�������Ŀ�������ω����/frh/gu�i/whitehome.png)�`g�yϋϝϯπ@�pointR����ϰ��+ߺ�  A�direc��g�yߋ�8�߯�>�/inQ��������0��E�choicQ�o��������@�touchup_�����+��=���@�arwrg��w���������F� ���� $6H�� l~����U� � 2D�hz �����c�
/ /./@/R/�v/�/�/ �/�/�/_/�/??*? <?N?`?7�e?�?�?�? �?�?�?�/
OO.O@O ROdO�?�O�O�O�O�O �OqO�O_*_<_N_`_ r__�_�_�_�_�_�_ _o&o8oJo\ono�_ �o�o�o�o�o�o�o�o "4FXj|� �������0� B�T�f�x�������� ҏ������,�>�P� b�t��������Ο�� �����:�L�^�p�h����/����:���ۯ�8�ɯ�(��7�,�S��POINT\���Ϫ����ο��  CHOI�CE]��TOUCHUP��8� \�Cπ�gϤ϶ϝ��� �������4��X�j��Qߎ�m;��whitehom^��������������poinf�R�d�v��� %������������� <�N�`�r�������7�>5�choic�������'*�4�t?ouchup��e�w���,�4�arwrgA��� /2�Sew�� �<���//+/ =/�a/s/�/�/�/�/ J/�/�/??'?9?�/ ]?o?�?�?�?�?�?X? �?�?O#O5OGO�?kO }O�O�O�O�O��bO�O __1_C_U_\Oy_�_ �_�_�_�_b_�_	oo -o?oQoco�_�o�o�o �o�o�opo); M_�o����� ��~�%�7�I�[� m��������Ǐُ� z��!�3�E�W�i�{� 
�����ß՟����� �/�A�S�e�w���� ����ѯ������+� =�O�a�s���������Ϳ߿�Ϟ��}������:�@L�^�6πϒ�l�,~� ��v��������A� (�e�w�^ߛ߂߿��� �������+��O�6� s�Z��������� ��O'�9�K�]�o��� �������������� ��5GYk}� ������1 CUgy��,� ���	//�?/Q/ c/u/�/�/(/�/�/�/ �/??)?�/M?_?q? �?�?�?6?�?�?�?O O%O�?IO[OmOO�O �O�ODO�O�O�O_!_ 3_�OW_i_{_�_�_�_ @_�_�_�_oo/oAo �eowo�o�o�o�o�_ �o�o+=O�o s�����\� ��'�9�K��o��� ������ɏۏj���� #�5�G�Y��}����� ��şןf�����1� C�U�g����������� ӯ�t�	��-�?�Q� c�򯇿������Ͽ� 󿂿�)�;�M�_�q�  ϕϧϹ�������~� �%�7�I�[�m��V`����V`����߼��ݦ������,��3���W�>�{� ��t���������� ��/�A�(�e�L����� ����������  =$asRo��� ��� �'9K ]o����� ���#/5/G/Y/k/ }//�/�/�/�/�/�/ ?�/1?C?U?g?y?�? ?�?�?�?�?�?	O�? -O?OQOcOuO�O�O(O �O�O�O�O__�O;_ M___q_�_�_$_�_�_ �_�_oo%o�_Io[o moo�o�o2o�o�o�o �o!�oEWi{ �������� �/�6S�e�w����� ����N������+� =�̏a�s��������� J�ߟ���'�9�K� ڟo���������ɯX� ����#�5�G�֯k� }�������ſ׿f��� ��1�C�U��yϋ� �ϯ�����b���	�� -�?�Q�c��χߙ߫� ������p���)�;� M�_��߃������h�����p����p����,�>��`�r�L�,^��V ����������!E W>{b���� ���/S: w�p����� //+/=/O/a/p�/ �/�/�/�/�/�/�/? '?9?K?]?o?�/�?�? �?�?�?�?|?O#O5O GOYOkO}OO�O�O�O �O�O�O�O_1_C_U_ g_y__�_�_�_�_�_ �_	o�_-o?oQocouo �oo�o�o�o�o�o �o);M_q�� $������� 7�I�[�m���� ��� Ǐُ����!��E� W�i�{�������ß՟ �����/���S�e� w�������<�ѯ��� ��+���O�a�s��� ������J�߿��� '�9�ȿ]�oρϓϥ� ��F��������#�5� G���k�}ߏߡ߳��� T�������1�C��� g�y��������b� ��	��-�?�Q���u� ����������^���@);M_6�a��6������������, ��7[mT �x�����/ !//E/,/i/{/b/�/ �/�/�/�/�/�/?? A?S?2�w?�?�?�?�? �?���?OO+O=OOO aO�?�O�O�O�O�O�O nO__'_9_K_]_�O �_�_�_�_�_�_�_|_ o#o5oGoYoko�_�o �o�o�o�o�oxo 1CUgy�� ������-�?� Q�c�u��������Ϗ �����)�;�M�_� q��������˟ݟ� ���%�7�I�[�m�� ��h?��ǯٯ���� �3�E�W�i�{����� .�ÿտ����Ϭ� A�S�e�wωϛ�*Ͽ� ��������+ߺ�O� a�s߅ߗߩ�8����� ����'��K�]�o� �����F������� �#�5���Y�k�}��� ����B������� 1C��gy��� �P��	-? �cu�����ڦ���������/-�@/R/,&,>?�/6?�/�/ �/�/�/?�/%?7?? [?B??�?x?�?�?�? �?�?O�?3OOWOiO PO�OtO�O�O���O�O __/_A_Pe_w_�_ �_�_�_�_`_�_oo +o=oOo�_so�o�o�o �o�o\o�o'9 K]�o����� �j��#�5�G�Y� �}�������ŏ׏� x���1�C�U�g��� ��������ӟ�t�	� �-�?�Q�c�u���� ����ϯ�󯂯�)� ;�M�_�q� ������� ˿ݿ���O%�7�I� [�m�φ��ϵ����� ����ߞ�3�E�W�i� {ߍ�߱��������� ��/�A�S�e�w�� ��*���������� ��=�O�a�s�����&� ��������'�� K]o���4� ���#�GY k}���B�� �//1/�U/g/y/ �/�/�/>/�/�/�/	?�?-???�A;�>����j?|? �=f?�?�?�6,�O�? �OO�?;OMO4OqOXO �O�O�O�O�O�O_�O %__I_[_B__f_�_ �_�_�_�_�_�_!o3o �Woio{o�o�o�o�/ �o�o�o/A�o ew����N� ���+�=��a�s� ��������͏\��� �'�9�K�ڏo����� ����ɟX�����#� 5�G�Y��}������� ůׯf�����1�C� U��y���������ӿ �t�	��-�?�Q�c� �ϙϫϽ�����p� ��)�;�M�_�q�Ho �ߧ߹���������� %�7�I�[�m���� �����������!�3� E�W�i�{�
������� ��������/AS ew����� ��+=Oas ��&����/ /�9/K/]/o/�/�/ "/�/�/�/�/�/?#? �/G?Y?k?}?�?�?0? �?�?�?�?OO�?CO�UOgOyO�O�O�O����K�������O�O�M�O _2_V,oc_o�_n_�_�_ �_�_�_oo�_;o"o _oqoXo�o|o�o�o�o �o�o�o7I0m T�������� �!�0OE�W�i�{��� ����@�Տ����� /���S�e�w������� <�џ�����+�=� ̟a�s���������J� ߯���'�9�ȯ]� o���������ɿX�� ���#�5�G�ֿk�}� �ϡϳ���T������ �1�C�U���yߋߝ� ������b���	��-� ?�Q���u����� ������)�;�M� _�f������������ ��~�%7I[m ��������z !3EWi{
 �������/ //A/S/e/w//�/�/ �/�/�/�/?�/+?=? O?a?s?�??�?�?�? �?�?O�?'O9OKO]O oO�O�O"O�O�O�O�O �O_�O5_G_Y_k_}_ �__�_�_�_�_�_o�o�$UI_IN�USER  ����@a��   o$o_�MENHIST �1D@e � ( M`���(/SOFTP�ART/GENL�INK?curr�ent=menu�page,153�,1_o�o�o�o�9)�o�o422�oU�gy�,xedi=t�bMAIND�8��� �'�/~71�[�m�����Q�o6�154J�������P��>�P�b� t�����'���Ο��� ����:�L�^�p��������4��a4�ѯ� ����+�.�O�a�s� ������8�Ϳ߿�� �'϶�ȿ]�oρϓ� �Ϸ�F��������#� 5���Y�k�}ߏߡ߳� B�T�������1�C� ��g�y�����אָ ����	��-�?�Q�T� u�����������^��� );M_��� �����l %7I[��� ����z/!/3/ E/W/i/��/�/�/�/ �/�/����?/?A?S? e?w?z/�?�?�?�?�? �?�?O+O=OOOaOsO �OO�O�O�O�O�O_ �O'_9_K_]_o_�__ �_�_�_�_�_�_o�_ 5oGoYoko}o�oo�o �o�o�o�o�/
?C Ugy���o�� ��	����Q�c� u�������:�Ϗ�� ��)���M�_�q��� ����6�H�ݟ��� %�7�Ɵ[�m������ ��D�ٯ����!�3����$UI_P�ANEDATA �1F���i��  	��}  frh/c�gtp/flex�dev.stm?�_width=0�&_height�=10����ice�=TP&_lin�es=15&_c�olumns=4���font=24�&_page=w�hole��E�!v)�  rim��  z�(�:�L�^�pς� 鿔ϸϟ����� �� ��6��Z�l�Sߐ�w����߭���!v� ��     ��"�}���J��2��39ཾ1ϵ/doub*�2���ual���$����� ����/���S�:�w� ��p����������� ��+OaH����
�   �i������ %xI��m� ���.���!/ /E/W/>/{/b/�/�/ �/�/�/�/�/?/?�I6k�fk?}?�?�? �?�??�?\OO1O COUOgO�?�O�O�O�O �O�O�O�O__?_&_ c_u_\_�_�_�_�_B? T?oo)o;oMo_o�_ �o�?�o�o�o�o�o zo7[B� x������� 3�E�,�i��_�_���� ÏՏ���L��/��o S�e�w��������џ ������+��O�a� H���l�������߯Ư �v���F�K�]�o��� ������ɿ<����� #�5�GϮ�k�}�dϡ� �����Ͼ������� C�U�<�y�`ߝ߯�"� 4�����	��-�?�� c�ֿ��������� ��Z����;�"�_�q� X���|�����������@%I�����T@������){ ��8J\n� �������/ �4//X/j/Q/�/u/��/�/�/�/x�������$UI_POST�YPE  ���� 	 ��/K?2QUICK�MEN  );�8?N?0RESTO�RE 1G���  ��*defaul�tx�DOUB�LE�=DUA�L�?medit�page,PART1,1�?*O<ONO|`OBmenuB154O�O�O�O�O �6�O�O__/_A_�1 �/R_d_�O�_�_�_�_ �_�_�_o/oAoSoeo o�o�o�o�o�o|_�o �oto=Oas� (������� '�9�K�]�o�|��� ���ۏ����#�Ə G�Y�k�}���2���ş ן��������,��� P�y���������d�� ��	��-�ЯQ�c�u�x����S=SCREi0�?n=u1�sc�0u2ڴ3�ڴ4ڴ5ڴ6ڴ7rڴ8ڱ��TAT%=�� }3��:UScER����Ӵksܳ�m�3m�4m�5m�6�m�7m�8m�0ND�O_CFG H�);d c0PD��W��Non�e\2N�_INFOW 1I���{00%���x�
�K�.� o߁�dߥ߷ߚ��߾� �����5�G�*�k�R<���OFFSET L)9�x�@��0 H�����������(� U�L�^���b������� ������$6��~?�p�
����_UFRAM�0@������RTOL_�ABRT���E�NB GRP �1M�9z1Cz  A�ec��cu ������h0�U/��MSK � 2�N��%���%Rs/ _'EVN2$�ƈ&v��2N��
 h���UEV!�td:\event_user\w/F� C7�/�B�F<��!SP�!�'sp�otweld=!C6????�0b$!b/�/�?�?�7!�? �?�?OAO�?�?wO"O �OFOXOjO�O�O_�O �O�OO_>_s__0_f_ �_�_�_�_�_o�_9o Ko�_o�o,o�oPobj~�&WRK 2OX�F�8�o	 �o @R-v�c�� �����*��N� `�;�����q���̏���ݏ���$VARS_CONFI���P�� FP@����CCRG��SP��Z@�9�D��B�BH�p����Ce���їϑ?�ᐶU�MRK2Y��)B�	��C�X��1: SC13?0EF2 *3�7��@����ch �5�B����A@��C�Ȑ� ��� ��9���ȯ�����"���ӑ��	�Z���� B��� u���z����᯾��� �Ϳ��*��'�`� ��Aϖρϓ������\�X�TCCc�ZR��4��pa��'�G�F,��![�� ��a 2345678901q�y�'9�n���n߰ߘ#����j�$����B��Ӗ ��ϑ?:�o=L{�� !p� �p��ia/[�� �Ԇ���������� )�;�(�:�q��p��� ���������%� I�[�H���{���������"�S�SELE�C�$!?�AVIoA_WO�`\T)�_ff,		��= �;G�P ��R'	�RTSYN'CSE�j��n�e�WINURL ?u��R����� //"�ISI�ONTMOU�/ ��*%c�]S۳��S۵@/� �FR:\,#\D�ATAs?MЄ� wMCk&LOGx/   UD1k&�EX�/��' ?B@ ���"�!�DESKTOP�-MC6FJ6K��/�#?%?�le �� n6  �����f�"�� -��N5K�   =���w1��t0� }�(TRAIN�/hH҆2�bd�3pw5>{4 #`�"'(:��^]� (���9 M��OO+O=OOO�O sO�O�O�O�O�O�O�O�_$(STAT _'� �z�b_t_�_�hq$�_�_'%_GES#�`]���0 �
����R�WHOMI}NV aS۾�`��b"���C�ז�&�WJMPERR� 2b]�
   =�jho^l��o�o�o �o�o�o�o.<�m`r�S_� R�EV cO^#�LEXr�Td7��1-e�_�VMPHASE � j���&�O�FFo_ENB � \�	P2R$e/SۿN��c|3�@:�`Q�u����?s33�4�1K� g�']g�t�g��&�S`�hWm�3�\BQ���C�F����81��_�
�A/�4��/�7k� B��C.�\@�4��� S�4�0�3��o�=�,������5ǟ[�s�C�;��Ԙ�#��rͫSAq��9��;�M�����Cj��ԓ�l��+&eB\�%�ՀS���_�u���������]�o��+��������%���6��+F�h_�����A�W������^Cr �B��+T�������*�dC�	Ml߯Կ�M�C�LA;B�6x��i敚,2��3��*ȹO��a�7�1�{�p������cda*�9�ӯɿ���C �����x�m�'�Y�K�	��e�Z����A�AC����Փ#�Ln��2A����Ϝ�����:6�B�������+�B)m�)�����C߀8�X��߄�� [��������3� ���i�^�p������ ������� /�!S� Hw�����y��� ���+=2a��_q��ÅTD�_FILTES`i��[ Է��P�� <//'/9/K/]/o/ �/�/�/6��/�/�/ ??,?>?P?b?t?�Y�SHIFTMENoU 1jWm<�|%��?�t�?�?O�? �?EOO.O{OROdO�O �O�O�O�O�O�O/__�	LIVE/S�NAP#Svsf�liv�~A_�^�PION &�U^PdRmenuz___��_�_�r�5G�kΉ�ֈ9MOG�l�~�z�łZDdm��a<�ۀ �P�$WA�ITDINEND�  �U��#bxfO9K-��oOUT�o�h�S�o�iTIM�e���lGo}�o2{��oz�oz�o�hREcLE�.��hTM^{�d�xc_ACT�WP-���h_DATA n΅�N�3�<E��RDIS�P�~��$XVRa�o9n�$ZABC_GRP 1p[k ,2J��=Qa��pVSPT q�9m���
�Z��_��Z)�?�އDCSCH`r#�����[IPbs[o!�۟���؊MPCF__G 1t����A0� O����u���Ġp�� 	�?���o`�  ?���2?�k��1�?�ɾ�����4/6��u��D5Oy���C���?����<� ���>%��6�����u=C������ί�1� ���	������˿� � 8��h�Ca���.~:��1�G�����۸��� &� �2�H�Vπ��,�>��0V�h��� �`�v����_CYLI�ND�w(� ��� ,(  * E�V��B��fߣߊ� ��������?� � ��D�+�=�z�ߞ�� ������g���@��'���v����̞�2x �� �=���? ��	��-=��`��zA��SPH�ERE 2y%�� ��*����X� kFX��|� ���///ew T/�x/_/q/�/��/��/�/��ZZ�v � f